module c499(sod0,sod1,sod2,sod3,sod4,sod5,sod6,sod7,sod8,sod9,sod10,sod11,sod12,sod13,sod14,sod15,sod16,sod17,sod18,sod19,sod20,sod21,sod22,sod23,sod24,sod25,sod26,sod27,sod28,sod29,sod30,sod31,sid0,sid1,sid2,sid3,sid4,sid5,sid6,sid7,sid8,sid9,sid10,sid11,sid12,sid13,sid14,sid15,sid16,sid17,sid18,sid19,sid20,sid21,sid22,sid23,sid24,sid25,sid26,sid27,sid28,sid29,sid30,sid31,sic0,sic1,sic2,sic3,sic4,sic5,sic6,sic7,sr);

  output sod0;
  output sod1;
  output sod2;
  output sod3;
  output sod4;
  output sod5;
  output sod6;
  output sod7;
  output sod8;
  output sod9;
  output sod10;
  output sod11;
  output sod12;
  output sod13;
  output sod14;
  output sod15;
  output sod16;
  output sod17;
  output sod18;
  output sod19;
  output sod20;
  output sod21;
  output sod22;
  output sod23;
  output sod24;
  output sod25;
  output sod26;
  output sod27;
  output sod28;
  output sod29;
  output sod30;
  output sod31;
  input sid0;
  input sid1;
  input sid2;
  input sid3;
  input sid4;
  input sid5;
  input sid6;
  input sid7;
  input sid8;
  input sid9;
  input sid10;
  input sid11;
  input sid12;
  input sid13;
  input sid14;
  input sid15;
  input sid16;
  input sid17;
  input sid18;
  input sid19;
  input sid20;
  input sid21;
  input sid22;
  input sid23;
  input sid24;
  input sid25;
  input sid26;
  input sid27;
  input sid28;
  input sid29;
  input sid30;
  input sid31;
  input sic0;
  input sic1;
  input sic2;
  input sic3;
  input sic4;
  input sic5;
  input sic6;
  input sic7;
  input sr;

  xor x0(sxa0,sid0,sid1);
  xor x1(sxa1,sid2,sid3);
  xor x2(sxa2,sid4,sid5);
  xor x3(sxa3,sid6,sid7);
  xor x4(sxa4,sid8,sid9);
  xor x5(sxa5,sid10,sid11);
  xor x6(sxa6,sid12,sid13);
  xor x7(sxa7,sid14,sid15);
  xor x8(sxa8,sid16,sid17);
  xor x9(sxa9,sid18,sid19);
  xor x10(sxa10,sid20,sid21);
  xor x11(sxa11,sid22,sid23);
  xor x12(sxa12,sid24,sid25);
  xor x13(sxa13,sid26,sid27);
  xor x14(sxa14,sid28,sid29);
  xor x15(sxa15,sid30,sid31);
  and x16(sh0,sic0,sr);
  and x17(sh1,sic1,sr);
  and x18(sh2,sic2,sr);
  and x19(sh3,sic3,sr);
  and x20(sh4,sic4,sr);
  and x21(sh5,sic5,sr);
  and x22(sh6,sic6,sr);
  and x23(sh7,sic7,sr);
  xor x24(sxb0,sid0,sid4);
  xor x25(sxc0,sid8,sid12);
  xor x26(sxb1,sid1,sid5);
  xor x27(sxc1,sid9,sid13);
  xor x28(sxb2,sid2,sid6);
  xor x29(sxc2,sid10,sid14);
  xor x30(sxb3,sid3,sid7);
  xor x31(sxc3,sid11,sid15);
  xor x32(sxb4,sid16,sid20);
  xor x33(sxc4,sid24,sid28);
  xor x34(sxb5,sid17,sid21);
  xor x35(sxc5,sid25,sid29);
  xor x36(sxb6,sid18,sid22);
  xor x37(sxc6,sid26,sid30);
  xor x38(sxb7,sid19,sid23);
  xor x39(sxc7,sid27,sid31);
  xor x40(sf0,sxa0,sxa1);
  xor x41(sf1,sxa2,sxa3);
  xor x42(sf2,sxa4,sxa5);
  xor x43(sf3,sxa6,sxa7);
  xor x44(sf4,sxa8,sxa9);
  xor x45(sf5,sxa10,sxa11);
  xor x46(sf6,sxa12,sxa13);
  xor x47(sf7,sxa14,sxa15);
  xor x48(sxe0,sxb0,sxc0);
  xor x49(sxe1,sxb1,sxc1);
  xor x50(sxe2,sxb2,sxc2);
  xor x51(sxe3,sxb3,sxc3);
  xor x52(sxe4,sxb4,sxc4);
  xor x53(sxe5,sxb5,sxc5);
  xor x54(sxe6,sxb6,sxc6);
  xor x55(sxe7,sxb7,sxc7);
  xor x56(sg0,sf0,sf1);
  xor x57(sg1,sf2,sf3);
  xor x58(sg2,sf0,sf2);
  xor x59(sg3,sf1,sf3);
  xor x60(sg4,sf4,sf5);
  xor x61(sg5,sf6,sf7);
  xor x62(sg6,sf4,sf6);
  xor x63(sg7,sf5,sf7);
  xor x64(sxd0,sh0,sg4);
  xor x65(sxd1,sh1,sg5);
  xor x66(sxd2,sh2,sg6);
  xor x67(sxd3,sh3,sg7);
  xor x68(sxd4,sh4,sg0);
  xor x69(sxd5,sh5,sg1);
  xor x70(sxd6,sh6,sg2);
  xor x71(sxd7,sh7,sg3);
  xor x72(ss0,sxe0,sxd0);
  xor x73(ss1,sxe1,sxd1);
  xor x74(ss2,sxe2,sxd2);
  xor x75(ss3,sxe3,sxd3);
  xor x76(ss4,sxe4,sxd4);
  xor x77(ss5,sxe5,sxd5);
  xor x78(ss6,sxe6,sxd6);
  xor x79(ss7,sxe7,sxd7);
  not x80(sy0a,ss0);
  not x81(sy1a,ss1);
  not x82(sy2a,ss2);
  not x83(sy0b,ss0);
  not x84(sy1b,ss1);
  not x85(sy3b,ss3);
  not x86(sy0c,ss0);
  not x87(sy2c,ss2);
  not x88(sy3c,ss3);
  not x89(sy1d,ss1);
  not x90(sy2d,ss2);
  not x91(sy3d,ss3);
  not x92(sy5i,ss5);
  not x93(sy7i,ss7);
  not x94(sy5j,ss5);
  not x95(sy6j,ss6);
  not x96(sy4k,ss4);
  not x97(sy7k,ss7);
  not x98(sy4l,ss4);
  not x99(sy6l,ss6);
  not x100(sy4a,ss4);
  not x101(sy5a,ss5);
  not x102(sy6a,ss6);
  not x103(sy4b,ss4);
  not x104(sy5b,ss5);
  not x105(sy7b,ss7);
  not x106(sy4c,ss4);
  not x107(sy6c,ss6);
  not x108(sy7c,ss7);
  not x109(sy5d,ss5);
  not x110(sy6d,ss6);
  not x111(sy7d,ss7);
  not x112(sy1i,ss1);
  not x113(sy3i,ss3);
  not x114(sy1j,ss1);
  not x115(sy2j,ss2);
  not x116(sy0k,ss0);
  not x117(sy3k,ss3);
  not x118(sy0l,ss0);
  not x119(sy2l,ss2);
  and x120(st0,sy0a,sy1a,sy2a,ss3);
  and x121(st1,sy0b,sy1b,ss2,sy3b);
  and x122(st2,sy0c,ss1,sy2c,sy3c);
  and x123(st3,ss0,sy1d,sy2d,sy3d);
  and x124(st4,sy4a,sy5a,sy6a,ss7);
  and x125(st5,sy4b,sy5b,ss6,sy7b);
  and x126(st6,sy4c,ss5,sy6c,sy7c);
  and x127(st7,ss4,sy5d,sy6d,sy7d);
  or x128(su0,st0,st1,st2,st3);
  or x129(su1,st4,st5,st6,st7);
  and x130(swa,ss4,sy5i,ss6,sy7i,su0);
  and x131(swb,ss4,sy5j,sy6j,ss7,su0);
  and x132(swc,sy4k,ss5,ss6,sy7k,su0);
  and x133(swd,sy4l,ss5,sy6l,ss7,su0);
  and x134(swe,ss0,sy1i,ss2,sy3i,su1);
  and x135(swf,ss0,sy1j,sy2j,ss3,su1);
  and x136(swg,sy0k,ss1,ss2,sy3k,su1);
  and x137(swh,sy0l,ss1,sy2l,ss3,su1);
  and x138(se0,ss0,swa);
  and x139(se1,ss1,swa);
  and x140(se2,ss2,swa);
  and x141(se3,ss3,swa);
  and x142(se4,ss0,swb);
  and x143(se5,ss1,swb);
  and x144(se6,ss2,swb);
  and x145(se7,ss3,swb);
  and x146(se8,ss0,swc);
  and x147(se9,ss1,swc);
  and x148(se10,ss2,swc);
  and x149(se11,ss3,swc);
  and x150(se12,ss0,swd);
  and x151(se13,ss1,swd);
  and x152(se14,ss2,swd);
  and x153(se15,ss3,swd);
  and x154(se16,ss4,swe);
  and x155(se17,ss5,swe);
  and x156(se18,ss6,swe);
  and x157(se19,ss7,swe);
  and x158(se20,ss4,swf);
  and x159(se21,ss5,swf);
  and x160(se22,ss6,swf);
  and x161(se23,ss7,swf);
  and x162(se24,ss4,swg);
  and x163(se25,ss5,swg);
  and x164(se26,ss6,swg);
  and x165(se27,ss7,swg);
  and x166(se28,ss4,swh);
  and x167(se29,ss5,swh);
  and x168(se30,ss6,swh);
  and x169(se31,ss7,swh);
  xor x170(sod0,sid0,se0);
  xor x171(sod1,sid1,se1);
  xor x172(sod2,sid2,se2);
  xor x173(sod3,sid3,se3);
  xor x174(sod4,sid4,se4);
  xor x175(sod5,sid5,se5);
  xor x176(sod6,sid6,se6);
  xor x177(sod7,sid7,se7);
  xor x178(sod8,sid8,se8);
  xor x179(sod9,sid9,se9);
  xor x180(sod10,sid10,se10);
  xor x181(sod11,sid11,se11);
  xor x182(sod12,sid12,se12);
  xor x183(sod13,sid13,se13);
  xor x184(sod14,sid14,se14);
  xor x185(sod15,sid15,se15);
  xor x186(sod16,sid16,se16);
  xor x187(sod17,sid17,se17);
  xor x188(sod18,sid18,se18);
  xor x189(sod19,sid19,se19);
  xor x190(sod20,sid20,se20);
  xor x191(sod21,sid21,se21);
  xor x192(sod22,sid22,se22);
  xor x193(sod23,sid23,se23);
  xor x194(sod24,sid24,se24);
  xor x195(sod25,sid25,se25);
  xor x196(sod26,sid26,se26);
  xor x197(sod27,sid27,se27);
  xor x198(sod28,sid28,se28);
  xor x199(sod29,sid29,se29);
  xor x200(sod30,sid30,se30);
  xor x201(sod31,sid31,se31);

endmodule
