module c2670(s169,s174,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s350,s335,s409,s369,s367,s411,s337,s384,s218,s219,s220,s221,s235,s236,s237,s238,s158,s259,s391,s173,s223,s234,s217,s325,s261,s319,s160,s162,s164,s166,s168,s171,s153,s176,s188,s299,s301,s286,s303,s288,s305,s290,s284,s321,s297,s280,s148,s282,s323,s156,s401,s227,s229,s311,s150,s145,s395,s295,s331,s397,s329,s231,s308,s225,s1,s2,s3,s4,s5,s6,s7,s8,s11,s14,s15,s16,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s32,s33,s34,s35,s36,s37,s40,s43,s44,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s60,s61,s62,s63,s64,s65,s66,s67,s68,s69,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s135,s136,s137,s138,s139,s140,s141,s142,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s452,s483,s543,s559,s567,s651,s661,s860,s868,s1083,s1341,s1348,s1384,s1956,s1961,s1966,s1971,s1976,s1981,s1986,s1991,s1996,s2066,s2067,s2072,s2078,s2084,s2090,s2096,s2100,s2104,s2105,s2106,s2427,s2430,s2435,s2438,s2443,s2446,s2451,s2454,s2474,s2678);

  inout s169;
  inout s174;
  output s177;
  output s178;
  output s179;
  output s180;
  output s181;
  output s182;
  output s183;
  output s184;
  output s185;
  output s186;
  output s189;
  output s190;
  output s191;
  output s192;
  output s193;
  output s194;
  output s195;
  output s196;
  output s197;
  output s198;
  output s199;
  output s200;
  output s201;
  output s202;
  output s203;
  output s204;
  output s205;
  output s206;
  output s207;
  output s208;
  output s209;
  output s210;
  output s211;
  output s212;
  output s213;
  output s214;
  output s215;
  output s239;
  output s240;
  output s241;
  output s242;
  output s243;
  output s244;
  output s245;
  output s246;
  output s247;
  output s248;
  output s249;
  output s250;
  output s251;
  output s252;
  output s253;
  output s254;
  output s255;
  output s256;
  output s257;
  output s262;
  output s263;
  output s264;
  output s265;
  output s266;
  output s267;
  output s268;
  output s269;
  output s270;
  output s271;
  output s272;
  output s273;
  output s274;
  output s275;
  output s276;
  output s277;
  output s278;
  output s279;
  output s350;
  output s335;
  output s409;
  output s369;
  output s367;
  output s411;
  output s337;
  output s384;
  output s218;
  output s219;
  output s220;
  output s221;
  output s235;
  output s236;
  output s237;
  output s238;
  output s158;
  output s259;
  output s391;
  output s173;
  output s223;
  output s234;
  output s217;
  output s325;
  output s261;
  output s319;
  output s160;
  output s162;
  output s164;
  output s166;
  output s168;
  output s171;
  output s153;
  output s176;
  output s188;
  output s299;
  output s301;
  output s286;
  output s303;
  output s288;
  output s305;
  output s290;
  output s284;
  output s321;
  output s297;
  output s280;
  output s148;
  output s282;
  output s323;
  output s156;
  output s401;
  output s227;
  output s229;
  output s311;
  output s150;
  output s145;
  output s395;
  output s295;
  output s331;
  output s397;
  output s329;
  output s231;
  output s308;
  output s225;
  input s1;
  input s2;
  input s3;
  input s4;
  input s5;
  input s6;
  input s7;
  input s8;
  input s11;
  input s14;
  input s15;
  input s16;
  input s19;
  input s20;
  input s21;
  input s22;
  input s23;
  input s24;
  input s25;
  input s26;
  input s27;
  input s28;
  input s29;
  input s32;
  input s33;
  input s34;
  input s35;
  input s36;
  input s37;
  input s40;
  input s43;
  input s44;
  input s47;
  input s48;
  input s49;
  input s50;
  input s51;
  input s52;
  input s53;
  input s54;
  input s55;
  input s56;
  input s57;
  input s60;
  input s61;
  input s62;
  input s63;
  input s64;
  input s65;
  input s66;
  input s67;
  input s68;
  input s69;
  input s72;
  input s73;
  input s74;
  input s75;
  input s76;
  input s77;
  input s78;
  input s79;
  input s80;
  input s81;
  input s82;
  input s85;
  input s86;
  input s87;
  input s88;
  input s89;
  input s90;
  input s91;
  input s92;
  input s93;
  input s94;
  input s95;
  input s96;
  input s99;
  input s100;
  input s101;
  input s102;
  input s103;
  input s104;
  input s105;
  input s106;
  input s107;
  input s108;
  input s111;
  input s112;
  input s113;
  input s114;
  input s115;
  input s116;
  input s117;
  input s118;
  input s119;
  input s120;
  input s123;
  input s124;
  input s125;
  input s126;
  input s127;
  input s128;
  input s129;
  input s130;
  input s131;
  input s132;
  input s135;
  input s136;
  input s137;
  input s138;
  input s139;
  input s140;
  input s141;
  input s142;
  input s177;
  input s178;
  input s179;
  input s180;
  input s181;
  input s182;
  input s183;
  input s184;
  input s185;
  input s186;
  input s189;
  input s190;
  input s191;
  input s192;
  input s193;
  input s194;
  input s195;
  input s196;
  input s197;
  input s198;
  input s199;
  input s200;
  input s201;
  input s202;
  input s203;
  input s204;
  input s205;
  input s206;
  input s207;
  input s208;
  input s209;
  input s210;
  input s211;
  input s212;
  input s213;
  input s214;
  input s215;
  input s239;
  input s240;
  input s241;
  input s242;
  input s243;
  input s244;
  input s245;
  input s246;
  input s247;
  input s248;
  input s249;
  input s250;
  input s251;
  input s252;
  input s253;
  input s254;
  input s255;
  input s256;
  input s257;
  input s262;
  input s263;
  input s264;
  input s265;
  input s266;
  input s267;
  input s268;
  input s269;
  input s270;
  input s271;
  input s272;
  input s273;
  input s274;
  input s275;
  input s276;
  input s277;
  input s278;
  input s279;
  input s452;
  input s483;
  input s543;
  input s559;
  input s567;
  input s651;
  input s661;
  input s860;
  input s868;
  input s1083;
  input s1341;
  input s1348;
  input s1384;
  input s1956;
  input s1961;
  input s1966;
  input s1971;
  input s1976;
  input s1981;
  input s1986;
  input s1991;
  input s1996;
  input s2066;
  input s2067;
  input s2072;
  input s2078;
  input s2084;
  input s2090;
  input s2096;
  input s2100;
  input s2104;
  input s2105;
  input s2106;
  input s2427;
  input s2430;
  input s2435;
  input s2438;
  input s2443;
  input s2446;
  input s2451;
  input s2454;
  input s2474;
  input s2678;

  buf x0(s350,s452);
  buf x1(s335,s452);
  buf x2(s409,s452);
  and x3(s546,s1,s3);
  not x4(s560,s559);
  buf x5(s369,s1083);
  buf x6(s367,s1083);
  not x7(s1385,s1384);
  buf x8(s411,s2066);
  buf x9(s337,s2066);
  buf x10(s384,s2066);
  and x11(s157,s2090,s2084,s2078,s2072);
  not x12(s547,s546);
  not x13(s218,s44);
  not x14(s219,s132);
  not x15(s220,s82);
  not x16(s221,s96);
  not x17(s235,s69);
  not x18(s236,s120);
  not x19(s237,s57);
  not x20(s238,s108);
  and x21(s258,s2,s15,s661);
  buf x22(s480,s661);
  and x23(s486,s37,s37);
  buf x24(s654,s452);
  buf x25(s655,s8);
  buf x26(s658,s8);
  buf x27(s772,s543);
  buf x28(s795,s651);
  not x29(s865,s860);
  not x30(s875,s868);
  and x31(s882,s11,s868);
  and x32(s1251,s132,s82,s96,s44);
  and x33(s1254,s120,s57,s108,s69);
  buf x34(s1261,s543);
  buf x35(s1284,s651);
  not x36(s1344,s1341);
  not x37(s1351,s1348);
  buf x38(s1394,s2104);
  buf x39(s1418,s2105);
  not x40(s2433,s2427);
  not x41(s2434,s2430);
  not x42(s2441,s2435);
  not x43(s2442,s2438);
  not x44(s2449,s2443);
  not x45(s2450,s2446);
  not x46(s2478,s2474);
  buf x47(s1631,s2104);
  buf x48(s1655,s2105);
  buf x49(s1710,s16);
  buf x50(s1721,s16);
  not x51(s2682,s2678);
  and x52(s1955,s7,s661);
  not x53(s1959,s1956);
  not x54(s1964,s1961);
  not x55(s1969,s1966);
  not x56(s1974,s1971);
  not x57(s1979,s1976);
  not x58(s1984,s1981);
  not x59(s1989,s1986);
  not x60(s1994,s1991);
  not x61(s1999,s1996);
  buf x62(s2001,s29);
  buf x63(s2012,s29);
  not x64(s2070,s2067);
  not x65(s2076,s2072);
  not x66(s2082,s2078);
  not x67(s2088,s2084);
  not x68(s2094,s2090);
  not x69(s2099,s2096);
  not x70(s2103,s2100);
  not x71(s2457,s2451);
  not x72(s2458,s2454);
  buf x73(s2461,s1348);
  buf x74(s2464,s1341);
  buf x75(s2471,s1956);
  buf x76(s2479,s1966);
  buf x77(s2482,s1961);
  buf x78(s2487,s1976);
  buf x79(s2490,s1971);
  buf x80(s2495,s1986);
  buf x81(s2498,s1981);
  buf x82(s2505,s1996);
  buf x83(s2508,s1991);
  buf x84(s2675,s2067);
  buf x85(s2683,s2078);
  buf x86(s2686,s2072);
  buf x87(s2691,s2090);
  buf x88(s2694,s2084);
  buf x89(s2699,s2100);
  buf x90(s2702,s2096);
  not x91(s158,s157);
  not x92(s259,s258);
  not x93(s487,s486);
  buf x94(s391,s654);
  nand x95(s1475,s2430,s2433);
  nand x96(s1476,s2427,s2434);
  nand x97(s1484,s2438,s2441);
  nand x98(s1485,s2435,s2442);
  nand x99(s1493,s2446,s2449);
  nand x100(s1494,s2443,s2450);
  nand x101(s2459,s2454,s2457);
  nand x102(s2460,s2451,s2458);
  and x103(s173,s94,s654);
  and x104(s216,s2106,s1955);
  not x105(s223,s1955);
  nand x106(s234,s567,s1955);
  not x107(s1253,s1251);
  not x108(s1256,s1254);
  and x109(s558,s1254,s1251);
  buf x110(s748,s655);
  not x111(s784,s772);
  not x112(s807,s795);
  and x113(s821,s80,s772,s795);
  and x114(s825,s68,s772,s795);
  and x115(s829,s79,s772,s795);
  and x116(s833,s78,s772,s795);
  and x117(s837,s77,s772,s795);
  and x118(s881,s11,s875);
  buf x119(s994,s655);
  not x120(s1273,s1261);
  not x121(s1296,s1284);
  and x122(s1310,s76,s1261,s1284);
  and x123(s1314,s75,s1261,s1284);
  and x124(s1318,s74,s1261,s1284);
  and x125(s1322,s73,s1261,s1284);
  and x126(s1326,s72,s1261,s1284);
  not x127(s1406,s1394);
  not x128(s1430,s1418);
  and x129(s1444,s114,s1394,s1418);
  and x130(s1448,s113,s1394,s1418);
  and x131(s1452,s112,s1394,s1418);
  and x132(s1456,s111,s1394,s1418);
  and x133(s1460,s1394,s1418);
  nand x134(s1477,s1475,s1476);
  nand x135(s1486,s1484,s1485);
  nand x136(s1495,s1493,s1494);
  not x137(s2477,s2471);
  nand x138(s1499,s2471,s2478);
  not x139(s2485,s2479);
  not x140(s2486,s2482);
  not x141(s2493,s2487);
  not x142(s2494,s2490);
  not x143(s1643,s1631);
  not x144(s1667,s1655);
  and x145(s1681,s118,s1631,s1655);
  and x146(s1685,s107,s1631,s1655);
  and x147(s1689,s117,s1631,s1655);
  and x148(s1693,s116,s1631,s1655);
  and x149(s1697,s115,s1631,s1655);
  not x150(s1716,s1710);
  not x151(s1728,s1721);
  not x152(s2681,s2675);
  nand x153(s1776,s2675,s2682);
  not x154(s2689,s2683);
  not x155(s2690,s2686);
  not x156(s2697,s2691);
  not x157(s2698,s2694);
  buf x158(s1831,s658);
  buf x159(s1893,s658);
  not x160(s2007,s2001);
  not x161(s2018,s2012);
  not x162(s2467,s2461);
  not x163(s2468,s2464);
  not x164(s2501,s2495);
  not x165(s2502,s2498);
  not x166(s2511,s2505);
  not x167(s2512,s2508);
  nand x168(s2518,s2459,s2460);
  buf x169(s2551,s1344);
  buf x170(s2559,s1351);
  buf x171(s2567,s1959);
  buf x172(s2575,s1964);
  buf x173(s2583,s1969);
  buf x174(s2591,s1974);
  buf x175(s2599,s1979);
  buf x176(s2607,s1984);
  buf x177(s2615,s1989);
  buf x178(s2623,s1994);
  not x179(s2705,s2699);
  not x180(s2706,s2702);
  buf x181(s2735,s1999);
  buf x182(s2743,s2070);
  buf x183(s2751,s2076);
  buf x184(s2759,s2082);
  buf x185(s2767,s2088);
  buf x186(s2775,s2094);
  not x187(s217,s216);
  and x188(s550,s2106,s1253);
  and x189(s552,s567,s1256);
  buf x190(s325,s558);
  or x191(s894,s881,s882);
  nand x192(s1498,s2474,s2477);
  nand x193(s1507,s2482,s2485);
  nand x194(s1508,s2479,s2486);
  nand x195(s1516,s2490,s2493);
  nand x196(s1517,s2487,s2494);
  nand x197(s1775,s2678,s2681);
  nand x198(s1784,s2686,s2689);
  nand x199(s1785,s2683,s2690);
  nand x200(s1793,s2694,s2697);
  nand x201(s1794,s2691,s2698);
  nand x202(s2469,s2464,s2467);
  nand x203(s2470,s2461,s2468);
  nand x204(s2503,s2498,s2501);
  nand x205(s2504,s2495,s2502);
  nand x206(s2513,s2508,s2511);
  nand x207(s2514,s2505,s2512);
  nand x208(s2707,s2702,s2705);
  nand x209(s2708,s2699,s2706);
  not x210(s261,s558);
  not x211(s551,s550);
  not x212(s553,s552);
  and x213(s818,s93,s784,s807);
  and x214(s819,s55,s772,s807);
  and x215(s820,s67,s784,s795);
  and x216(s822,s81,s784,s807);
  and x217(s823,s43,s772,s807);
  and x218(s824,s56,s784,s795);
  and x219(s826,s92,s784,s807);
  and x220(s827,s54,s772,s807);
  and x221(s828,s66,s784,s795);
  and x222(s830,s91,s784,s807);
  and x223(s831,s53,s772,s807);
  and x224(s832,s65,s784,s795);
  and x225(s834,s90,s784,s807);
  and x226(s835,s52,s772,s807);
  and x227(s836,s64,s784,s795);
  and x228(s1307,s89,s1273,s1296);
  and x229(s1308,s51,s1261,s1296);
  and x230(s1309,s63,s1273,s1284);
  and x231(s1311,s88,s1273,s1296);
  and x232(s1312,s50,s1261,s1296);
  and x233(s1313,s62,s1273,s1284);
  and x234(s1315,s87,s1273,s1296);
  and x235(s1316,s49,s1261,s1296);
  and x236(s1317,s1273,s1284);
  and x237(s1319,s86,s1273,s1296);
  and x238(s1320,s48,s1261,s1296);
  and x239(s1321,s61,s1273,s1284);
  and x240(s1323,s85,s1273,s1296);
  and x241(s1324,s47,s1261,s1296);
  and x242(s1325,s60,s1273,s1284);
  and x243(s1441,s138,s1406,s1430);
  and x244(s1442,s102,s1394,s1430);
  and x245(s1443,s126,s1406,s1418);
  and x246(s1445,s137,s1406,s1430);
  and x247(s1446,s101,s1394,s1430);
  and x248(s1447,s125,s1406,s1418);
  and x249(s1449,s136,s1406,s1430);
  and x250(s1450,s100,s1394,s1430);
  and x251(s1451,s124,s1406,s1418);
  and x252(s1453,s135,s1406,s1430);
  and x253(s1454,s99,s1394,s1430);
  and x254(s1455,s123,s1406,s1418);
  and x255(s1457,s1406,s1430);
  and x256(s1458,s1394,s1430);
  and x257(s1459,s1406,s1418);
  not x258(s1481,s1477);
  not x259(s1490,s1486);
  nand x260(s1500,s1498,s1499);
  nand x261(s1509,s1507,s1508);
  nand x262(s1518,s1516,s1517);
  buf x263(s1521,s1495);
  buf x264(s1525,s1495);
  not x265(s2557,s2551);
  not x266(s2565,s2559);
  not x267(s2573,s2567);
  not x268(s2581,s2575);
  not x269(s2589,s2583);
  not x270(s2597,s2591);
  not x271(s2605,s2599);
  not x272(s2613,s2607);
  not x273(s2621,s2615);
  not x274(s2629,s2623);
  and x275(s1678,s142,s1643,s1667);
  and x276(s1679,s106,s1631,s1667);
  and x277(s1680,s130,s1643,s1655);
  and x278(s1682,s131,s1643,s1667);
  and x279(s1683,s95,s1631,s1667);
  and x280(s1684,s119,s1643,s1655);
  and x281(s1686,s141,s1643,s1667);
  and x282(s1687,s105,s1631,s1667);
  and x283(s1688,s129,s1643,s1655);
  and x284(s1690,s140,s1643,s1667);
  and x285(s1691,s104,s1631,s1667);
  and x286(s1692,s128,s1643,s1655);
  and x287(s1694,s139,s1643,s1667);
  and x288(s1695,s103,s1631,s1667);
  and x289(s1696,s127,s1643,s1655);
  and x290(s1734,s19,s1716);
  and x291(s1736,s4,s1716);
  and x292(s1738,s20,s1716);
  and x293(s1740,s5,s1716);
  and x294(s1742,s21,s1728);
  and x295(s1744,s22,s1728);
  and x296(s1746,s23,s1728);
  and x297(s1748,s6,s1728);
  and x298(s1750,s24,s1728);
  nand x299(s1777,s1775,s1776);
  nand x300(s1786,s1784,s1785);
  nand x301(s1795,s1793,s1794);
  and x302(s2023,s25,s2007);
  and x303(s2025,s32,s2007);
  and x304(s2027,s26,s2007);
  and x305(s2029,s33,s2007);
  and x306(s2031,s27,s2018);
  and x307(s2033,s34,s2018);
  and x308(s2035,s35,s2018);
  and x309(s2037,s28,s2018);
  not x310(s2741,s2735);
  not x311(s2749,s2743);
  not x312(s2757,s2751);
  not x313(s2765,s2759);
  not x314(s2773,s2767);
  not x315(s2781,s2775);
  nand x316(s2515,s2469,s2470);
  not x317(s2522,s2518);
  nand x318(s2525,s2513,s2514);
  nand x319(s2528,s2503,s2504);
  nand x320(s2730,s2707,s2708);
  and x321(s554,s551,s553);
  or x322(s838,s818,s819,s820,s821);
  or x323(s841,s822,s823,s824,s825);
  or x324(s846,s826,s827,s828,s829);
  or x325(s854,s830,s831,s832,s833);
  or x326(s857,s834,s835,s836,s837);
  or x327(s1327,s1307,s1308,s1309,s1310);
  or x328(s1329,s1311,s1312,s1313,s1314);
  or x329(s1331,s1315,s1316,s1317,s1318);
  or x330(s1333,s1319,s1320,s1321,s1322);
  or x331(s1335,s1323,s1324,s1325,s1326);
  or x332(s1461,s1441,s1442,s1443,s1444);
  or x333(s1464,s1445,s1446,s1447,s1448);
  or x334(s1467,s1449,s1450,s1451,s1452);
  or x335(s1470,s1453,s1454,s1455,s1456);
  or x336(s1473,s1457,s1458,s1459,s1460);
  or x337(s1698,s1682,s1683,s1684,s1685);
  or x338(s1701,s1686,s1687,s1688,s1689);
  or x339(s1704,s1690,s1691,s1692,s1693);
  or x340(s1707,s1694,s1695,s1696,s1697);
  or x341(s2634,s1678,s1679,s1680,s1681);
  buf x342(s319,s554);
  not x343(s1504,s1500);
  not x344(s1513,s1509);
  not x345(s1524,s1521);
  not x346(s1528,s1525);
  buf x347(s1529,s1518);
  buf x348(s1533,s1518);
  and x349(s1538,s1486,s1477,s1521);
  and x350(s1541,s1490,s1481,s1525);
  not x351(s1781,s1777);
  not x352(s1790,s1786);
  buf x353(s1806,s1795);
  buf x354(s1810,s1795);
  not x355(s2734,s2730);
  not x356(s2521,s2515);
  nand x357(s2524,s2515,s2522);
  not x358(s2531,s2525);
  not x359(s2532,s2528);
  and x360(s144,s838,s860);
  and x361(s147,s846,s860);
  and x362(s152,s841,s860);
  not x363(s160,s1464);
  not x364(s162,s1467);
  not x365(s164,s1461);
  not x366(s166,s1329);
  not x367(s168,s1327);
  not x368(s171,s857);
  and x369(s175,s480,s483,s36,s554);
  and x370(s187,s480,s483,s554,s547);
  buf x371(s516,s838);
  not x372(s852,s846);
  and x373(s885,s841,s875);
  and x374(s887,s846,s875);
  and x375(s893,s1327,s868);
  not x376(s1028,s838);
  not x377(s1031,s841);
  not x378(s1035,s846);
  buf x379(s1041,s854);
  buf x380(s1049,s857);
  buf x381(s1057,s1327);
  buf x382(s1060,s1329);
  buf x383(s1066,s1331);
  buf x384(s1072,s1333);
  buf x385(s1078,s1335);
  nand x386(s1213,s2099,s1470);
  nand x387(s1218,s2103,s1473);
  buf x388(s1250,s1704);
  and x389(s1387,s1461,s1385);
  not x390(s1389,s1464);
  and x391(s1537,s1481,s1486,s1524);
  and x392(s1540,s1477,s1490,s1528);
  and x393(s1735,s841,s1710);
  and x394(s1737,s846,s1710);
  and x395(s1739,s854,s1710);
  and x396(s1741,s857,s1710);
  and x397(s1743,s1327,s1721);
  and x398(s1745,s1329,s1721);
  and x399(s1747,s1331,s1721);
  and x400(s1749,s1333,s1721);
  and x401(s1751,s1335,s1721);
  not x402(s2638,s2634);
  and x403(s2024,s1698,s2001);
  and x404(s2026,s1701,s2001);
  and x405(s2028,s1704,s2001);
  and x406(s2030,s1707,s2001);
  and x407(s2032,s1461,s2012);
  and x408(s2034,s1464,s2012);
  and x409(s2036,s1467,s2012);
  and x410(s2038,s1470,s2012);
  buf x411(s2154,s841);
  nand x412(s2523,s2518,s2521);
  nand x413(s2533,s2528,s2531);
  nand x414(s2534,s2525,s2532);
  buf x415(s2631,s1698);
  buf x416(s2639,s1704);
  buf x417(s2642,s1701);
  buf x418(s2647,s1461);
  buf x419(s2650,s1707);
  buf x420(s2655,s1467);
  buf x421(s2658,s1464);
  buf x422(s2665,s1473);
  buf x423(s2668,s1470);
  or x424(s153,s865,s152);
  not x425(s176,s175);
  not x426(s188,s187);
  buf x427(s299,s1041);
  buf x428(s301,s1049);
  buf x429(s286,s1057);
  buf x430(s303,s1060);
  buf x431(s288,s1066);
  buf x432(s305,s1072);
  buf x433(s290,s1078);
  not x434(s1532,s1529);
  not x435(s1536,s1533);
  nor x436(s1539,s1537,s1538);
  nor x437(s1542,s1540,s1541);
  and x438(s1544,s1509,s1500,s1529);
  and x439(s1547,s1513,s1504,s1533);
  or x440(s2065,s2037,s2038);
  not x441(s1809,s1806);
  not x442(s1813,s1810);
  and x443(s1821,s1786,s1777,s1806);
  and x444(s1824,s1790,s1781,s1810);
  nand x445(s2538,s2523,s2524);
  nand x446(s2546,s2533,s2534);
  or x447(s2554,s1734,s1735);
  or x448(s2562,s1736,s1737);
  or x449(s2570,s1738,s1739);
  or x450(s2578,s1740,s1741);
  or x451(s2586,s1742,s1743);
  or x452(s2594,s1744,s1745);
  or x453(s2602,s1746,s1747);
  or x454(s2610,s1748,s1749);
  or x455(s2618,s1750,s1751);
  or x456(s2626,s2023,s2024);
  or x457(s2738,s2025,s2026);
  or x458(s2746,s2027,s2028);
  or x459(s2754,s2029,s2030);
  or x460(s2762,s2031,s2032);
  or x461(s2770,s2033,s2034);
  or x462(s2778,s2035,s2036);
  and x463(s456,s1389,s1387,s40);
  not x464(s466,s1387);
  nand x465(s562,s560,s852);
  and x466(s883,s516,s875);
  and x467(s889,s1049,s868);
  and x468(s891,s1041,s875);
  not x469(s1043,s1041);
  not x470(s1051,s1049);
  not x471(s1062,s1060);
  not x472(s1068,s1066);
  not x473(s1074,s1072);
  not x474(s1080,s1078);
  and x475(s1225,s2099,s1213);
  and x476(s1227,s1213,s1470);
  and x477(s1232,s2103,s1218);
  and x478(s1234,s1218,s1473);
  and x479(s1543,s1504,s1509,s1532);
  and x480(s1546,s1500,s1513,s1536);
  not x481(s2637,s2631);
  nand x482(s1753,s2631,s2638);
  not x483(s2645,s2639);
  not x484(s2646,s2642);
  not x485(s2653,s2647);
  not x486(s2654,s2650);
  and x487(s1820,s1781,s1786,s1809);
  and x488(s1823,s1777,s1790,s1813);
  buf x489(s2107,s1031);
  buf x490(s2110,s1028);
  buf x491(s2118,s1035);
  not x492(s2123,s1057);
  not x493(s2151,s852);
  not x494(s2158,s2154);
  buf x495(s2161,s1031);
  buf x496(s2164,s1028);
  buf x497(s2172,s1035);
  buf x498(s2235,s516);
  buf x499(s2262,s1035);
  buf x500(s2350,s1035);
  nand x501(s2535,s1542,s1539);
  not x502(s2661,s2655);
  not x503(s2662,s2658);
  not x504(s2671,s2665);
  not x505(s2672,s2668);
  and x506(s468,s40,s1389,s466);
  or x507(s897,s887,s889);
  or x508(s898,s891,s893);
  or x509(s1228,s1225,s1227);
  or x510(s1235,s1232,s1234);
  nor x511(s1545,s1543,s1544);
  nor x512(s1548,s1546,s1547);
  not x513(s2542,s2538);
  not x514(s2550,s2546);
  nand x515(s1561,s2554,s2557);
  not x516(s2558,s2554);
  nand x517(s1565,s2562,s2565);
  not x518(s2566,s2562);
  nand x519(s1569,s2570,s2573);
  not x520(s2574,s2570);
  nand x521(s1573,s2578,s2581);
  not x522(s2582,s2578);
  nand x523(s1577,s2586,s2589);
  not x524(s2590,s2586);
  nand x525(s1581,s2594,s2597);
  not x526(s2598,s2594);
  nand x527(s1585,s2602,s2605);
  not x528(s2606,s2602);
  nand x529(s1589,s2610,s2613);
  not x530(s2614,s2610);
  nand x531(s1593,s2618,s2621);
  not x532(s2622,s2618);
  nand x533(s1597,s2626,s2629);
  not x534(s2630,s2626);
  nand x535(s1752,s2634,s2637);
  nand x536(s1761,s2642,s2645);
  nand x537(s1762,s2639,s2646);
  nand x538(s1770,s2650,s2653);
  nand x539(s1771,s2647,s2654);
  nor x540(s1822,s1820,s1821);
  nor x541(s1825,s1823,s1824);
  nand x542(s2039,s2738,s2741);
  not x543(s2742,s2738);
  nand x544(s2043,s2746,s2749);
  not x545(s2750,s2746);
  nand x546(s2047,s2754,s2757);
  not x547(s2758,s2754);
  nand x548(s2051,s2762,s2765);
  not x549(s2766,s2762);
  nand x550(s2055,s2770,s2773);
  not x551(s2774,s2770);
  nand x552(s2059,s2778,s2781);
  not x553(s2782,s2778);
  nand x554(s2663,s2658,s2661);
  nand x555(s2664,s2655,s2662);
  nand x556(s2673,s2668,s2671);
  nand x557(s2674,s2665,s2672);
  and x558(s146,s562,s865);
  not x559(s462,s456);
  not x560(s2113,s2107);
  not x561(s2114,s2110);
  not x562(s2122,s2118);
  not x563(s2129,s2123);
  buf x564(s592,s562);
  not x565(s2167,s2161);
  not x566(s2168,s2164);
  not x567(s2176,s2172);
  not x568(s2241,s2235);
  not x569(s2266,s2262);
  not x570(s743,s456);
  buf x571(s749,s456);
  and x572(s886,s562,s868);
  buf x573(s284,s897);
  buf x574(s321,s897);
  buf x575(s297,s898);
  buf x576(s280,s898);
  buf x577(s995,s456);
  not x578(s1006,s456);
  nand x579(s1550,s2535,s2542);
  not x580(s2354,s2350);
  not x581(s2541,s2535);
  nand x582(s1562,s2551,s2558);
  nand x583(s1566,s2559,s2566);
  nand x584(s1570,s2567,s2574);
  nand x585(s1574,s2575,s2582);
  nand x586(s1578,s2583,s2590);
  nand x587(s1582,s2591,s2598);
  nand x588(s1586,s2599,s2606);
  nand x589(s1590,s2607,s2614);
  nand x590(s1594,s2615,s2622);
  nand x591(s1598,s2623,s2630);
  nand x592(s1754,s1752,s1753);
  nand x593(s1763,s1761,s1762);
  nand x594(s1772,s1770,s1771);
  nand x595(s2040,s2735,s2742);
  nand x596(s2044,s2743,s2750);
  nand x597(s2048,s2751,s2758);
  nand x598(s2052,s2759,s2766);
  nand x599(s2056,s2767,s2774);
  nand x600(s2060,s2775,s2782);
  buf x601(s2115,s1043);
  buf x602(s2126,s1051);
  buf x603(s2131,s1068);
  buf x604(s2134,s1062);
  buf x605(s2141,s1080);
  buf x606(s2144,s1074);
  not x607(s2157,s2151);
  nand x608(s2160,s2151,s2158);
  buf x609(s2169,s1043);
  buf x610(s2177,s1068);
  buf x611(s2180,s1062);
  buf x612(s2187,s1080);
  buf x613(s2190,s1074);
  not x614(s2207,s562);
  buf x615(s2254,s1043);
  buf x616(s2334,s1051);
  buf x617(s2342,s1043);
  buf x618(s2422,s1051);
  nand x619(s2543,s1548,s1545);
  nand x620(s2709,s2673,s2674);
  nand x621(s2712,s2663,s2664);
  nand x622(s2727,s1825,s1822);
  or x623(s148,s146,s147);
  nand x624(s569,s2110,s2113);
  nand x625(s570,s2107,s2114);
  nand x626(s599,s2164,s2167);
  nand x627(s600,s2161,s2168);
  or x628(s896,s885,s886);
  nand x629(s1549,s2538,s2541);
  not x630(s1243,s1228);
  not x631(s1245,s1235);
  buf x632(s1257,s468);
  buf x633(s1258,s468);
  nand x634(s1563,s1561,s1562);
  nand x635(s1567,s1565,s1566);
  nand x636(s1571,s1569,s1570);
  nand x637(s1575,s1573,s1574);
  nand x638(s1579,s1577,s1578);
  nand x639(s1583,s1581,s1582);
  nand x640(s1587,s1585,s1586);
  nand x641(s1591,s1589,s1590);
  nand x642(s1595,s1593,s1594);
  nand x643(s1599,s1597,s1598);
  nand x644(s2041,s2039,s2040);
  nand x645(s2045,s2043,s2044);
  nand x646(s2049,s2047,s2048);
  nand x647(s2053,s2051,s2052);
  nand x648(s2057,s2055,s2056);
  nand x649(s2061,s2059,s2060);
  nand x650(s2159,s2154,s2157);
  buf x651(s475,s462);
  and x652(s490,s1078,s743);
  and x653(s496,s1698,s743);
  and x654(s502,s1701,s743);
  and x655(s508,s1250,s743);
  and x656(s765,s1057,s749);
  and x657(s769,s1060,s749);
  nand x658(s571,s569,s570);
  not x659(s2121,s2115);
  nand x660(s579,s2115,s2122);
  nand x661(s587,s2126,s2129);
  not x662(s2130,s2126);
  not x663(s596,s592);
  nand x664(s601,s599,s600);
  not x665(s2175,s2169);
  nand x666(s609,s2169,s2176);
  not x667(s2258,s2254);
  and x668(s1014,s1057,s995);
  and x669(s1018,s1060,s995);
  and x670(s717,s1078,s1006);
  and x671(s723,s1698,s1006);
  and x672(s729,s1701,s1006);
  and x673(s735,s1250,s1006);
  not x674(s753,s749);
  buf x675(s282,s896);
  buf x676(s323,s896);
  not x677(s2338,s2334);
  not x678(s999,s995);
  nand x679(s1091,s1549,s1550);
  not x680(s2346,s2342);
  not x681(s2426,s2422);
  buf x682(s1337,s462);
  not x683(s2549,s2543);
  nand x684(s1552,s2543,s2550);
  not x685(s1600,s1599);
  not x686(s1596,s1595);
  not x687(s1592,s1591);
  not x688(s1588,s1587);
  not x689(s1584,s1583);
  not x690(s1580,s1579);
  not x691(s1576,s1575);
  not x692(s1572,s1571);
  not x693(s1568,s1567);
  not x694(s1564,s1563);
  not x695(s2062,s2061);
  not x696(s2058,s2057);
  not x697(s2054,s2053);
  not x698(s2050,s2049);
  not x699(s2046,s2045);
  not x700(s2042,s2041);
  not x701(s1758,s1754);
  not x702(s1767,s1763);
  buf x703(s1798,s1772);
  buf x704(s1802,s1772);
  not x705(s2733,s2727);
  nand x706(s1829,s2727,s2734);
  not x707(s2137,s2131);
  not x708(s2138,s2134);
  not x709(s2147,s2141);
  not x710(s2148,s2144);
  not x711(s2183,s2177);
  not x712(s2184,s2180);
  not x713(s2193,s2187);
  not x714(s2194,s2190);
  nand x715(s2210,s2159,s2160);
  not x716(s2213,s2207);
  not x717(s2715,s2709);
  not x718(s2716,s2712);
  and x719(s1094,s1235,s1245);
  and x720(s1096,s1228,s1243);
  nand x721(s578,s2118,s2121);
  nand x722(s588,s2123,s2130);
  nand x723(s608,s2172,s2175);
  buf x724(s742,s1257);
  buf x725(s1005,s1257);
  not x726(s1092,s1091);
  nand x727(s1551,s2546,s2549);
  and x728(s1554,s1600,s1596,s1592,s1588,s1584);
  and x729(s1555,s1580,s1576,s1572,s1568,s1564);
  and x730(s1557,s2065,s2062);
  and x731(s1558,s2058,s2054,s2050,s2046,s2042);
  nand x732(s1828,s2730,s2733);
  buf x733(s1845,s1258);
  buf x734(s1907,s1258);
  nand x735(s2139,s2134,s2137);
  nand x736(s2140,s2131,s2138);
  nand x737(s2149,s2144,s2147);
  nand x738(s2150,s2141,s2148);
  nand x739(s2185,s2180,s2183);
  nand x740(s2186,s2177,s2184);
  nand x741(s2195,s2190,s2193);
  nand x742(s2196,s2187,s2194);
  nand x743(s2717,s2712,s2715);
  nand x744(s2718,s2709,s2716);
  or x745(s154,s1094,s1245);
  or x746(s155,s1096,s1243);
  and x747(s763,s1057,s753);
  and x748(s767,s1060,s753);
  and x749(s531,s1066,s753);
  and x750(s537,s1072,s753);
  not x751(s575,s571);
  nand x752(s580,s578,s579);
  nand x753(s589,s587,s588);
  not x754(s605,s601);
  nand x755(s610,s608,s609);
  and x756(s1012,s1057,s999);
  and x757(s1016,s1060,s999);
  and x758(s705,s1066,s999);
  and x759(s711,s1072,s999);
  and x760(s1093,s1092,s14);
  buf x761(s1355,s475);
  nand x762(s1553,s1551,s1552);
  and x763(s1556,s1554,s1555);
  and x764(s1559,s1557,s1558);
  buf x765(s1601,s1337);
  not x766(s1801,s1798);
  not x767(s1805,s1802);
  and x768(s1815,s1763,s1754,s1798);
  and x769(s1818,s1767,s1758,s1802);
  nand x770(s1830,s1828,s1829);
  buf x771(s1836,s475);
  buf x772(s1850,s475);
  buf x773(s1898,s1337);
  buf x774(s1912,s1337);
  nand x775(s2197,s2149,s2150);
  nand x776(s2200,s2139,s2140);
  not x777(s2214,s2210);
  nand x778(s2215,s2210,s2213);
  nand x779(s2217,s2195,s2196);
  nand x780(s2220,s2185,s2186);
  nand x781(s2722,s2717,s2718);
  nand x782(s156,s154,s155);
  and x783(s492,s490,s742);
  and x784(s498,s496,s742);
  and x785(s504,s502,s742);
  and x786(s510,s508,s742);
  or x787(s519,s763,s765);
  or x788(s525,s767,s769);
  and x789(s533,s531,s748);
  and x790(s539,s537,s748);
  or x791(s693,s1012,s1014);
  or x792(s699,s1016,s1018);
  and x793(s707,s705,s994);
  and x794(s713,s711,s994);
  and x795(s719,s717,s1005);
  and x796(s725,s723,s1005);
  and x797(s731,s729,s1005);
  and x798(s737,s735,s1005);
  buf x799(s401,s1093);
  and x800(s1560,s1556,s1559,s894);
  and x801(s1814,s1758,s1763,s1801);
  and x802(s1817,s1754,s1767,s1805);
  nand x803(s2216,s2207,s2214);
  not x804(s227,s1830);
  not x805(s229,s1553);
  not x806(s493,s492);
  not x807(s499,s498);
  not x808(s505,s504);
  not x809(s511,s510);
  and x810(s521,s519,s748);
  and x811(s527,s525,s748);
  not x812(s534,s533);
  not x813(s540,s539);
  not x814(s584,s580);
  buf x815(s613,s589);
  buf x816(s617,s589);
  buf x817(s621,s610);
  buf x818(s625,s610);
  and x819(s676,s1344,s1355);
  and x820(s695,s693,s994);
  and x821(s701,s699,s994);
  not x822(s708,s707);
  not x823(s714,s713);
  not x824(s720,s719);
  not x825(s726,s725);
  not x826(s732,s731);
  not x827(s738,s737);
  not x828(s1087,s1093);
  and x829(s1108,s1344,s1601);
  not x830(s1361,s1355);
  and x831(s1369,s1351,s1355);
  and x832(s1373,s1959,s1355);
  and x833(s1377,s1964,s1355);
  buf x834(s311,s1560);
  not x835(s1607,s1601);
  and x836(s1615,s1351,s1601);
  and x837(s1619,s1959,s1601);
  and x838(s1623,s1964,s1601);
  nor x839(s1816,s1814,s1815);
  nor x840(s1819,s1817,s1818);
  not x841(s2726,s2722);
  not x842(s1842,s1836);
  and x843(s1858,s1969,s1836);
  and x844(s1863,s1974,s1836);
  and x845(s1866,s1979,s1836);
  and x846(s1868,s1984,s1836);
  and x847(s1870,s1989,s1850);
  and x848(s1872,s1994,s1850);
  and x849(s1874,s1999,s1850);
  and x850(s1876,s2070,s1850);
  not x851(s1904,s1898);
  and x852(s1920,s1969,s1898);
  and x853(s1925,s1974,s1898);
  and x854(s1928,s1979,s1898);
  and x855(s1930,s1984,s1898);
  and x856(s1932,s1989,s1912);
  and x857(s1934,s1994,s1912);
  and x858(s1936,s1999,s1912);
  and x859(s1938,s2070,s1912);
  not x860(s2203,s2197);
  not x861(s2204,s2200);
  not x862(s2223,s2217);
  not x863(s2224,s2220);
  nand x864(s2238,s2215,s2216);
  not x865(s150,s1560);
  not x866(s522,s521);
  not x867(s528,s527);
  not x868(s696,s695);
  not x869(s702,s701);
  and x870(s1881,s1866,s1831);
  and x871(s1883,s1868,s1831);
  and x872(s1885,s1870,s1845);
  and x873(s1887,s1872,s1845);
  and x874(s1889,s1874,s1845);
  and x875(s1891,s1876,s1845);
  and x876(s1943,s1928,s1893);
  and x877(s1945,s1930,s1893);
  and x878(s1947,s1932,s1907);
  and x879(s1949,s1934,s1907);
  and x880(s1951,s1936,s1907);
  and x881(s1953,s1938,s1907);
  nand x882(s2205,s2200,s2203);
  nand x883(s2206,s2197,s2204);
  nand x884(s2225,s2220,s2223);
  nand x885(s2226,s2217,s2224);
  nand x886(s2719,s1819,s1816);
  not x887(s616,s613);
  not x888(s620,s617);
  not x889(s624,s621);
  not x890(s628,s625);
  and x891(s630,s580,s571,s613);
  and x892(s633,s584,s575,s617);
  and x893(s636,s601,s592,s621);
  and x894(s639,s605,s596,s625);
  nand x895(s645,s2238,s2241);
  not x896(s2242,s2238);
  and x897(s675,s1999,s1361);
  and x898(s1107,s1999,s1607);
  and x899(s1368,s2070,s1361);
  and x900(s1371,s2076,s1361);
  and x901(s1375,s2082,s1361);
  and x902(s1614,s2070,s1607);
  and x903(s1617,s2076,s1607);
  and x904(s1621,s2082,s1607);
  and x905(s1856,s2088,s1842);
  and x906(s1861,s2094,s1842);
  and x907(s1918,s2088,s1904);
  and x908(s1923,s2094,s1904);
  nand x909(s2230,s2205,s2206);
  nand x910(s2246,s2225,s2226);
  buf x911(s2270,s511);
  buf x912(s2278,s505);
  buf x913(s2286,s499);
  buf x914(s2294,s493);
  buf x915(s2302,s540);
  buf x916(s2310,s534);
  buf x917(s2358,s738);
  buf x918(s2366,s732);
  buf x919(s2374,s726);
  buf x920(s2382,s720);
  buf x921(s2390,s714);
  buf x922(s2398,s708);
  and x923(s629,s575,s580,s616);
  and x924(s632,s571,s584,s620);
  and x925(s635,s596,s601,s624);
  and x926(s638,s592,s605,s628);
  nand x927(s646,s2235,s2242);
  or x928(s677,s675,s676);
  nand x929(s1827,s2719,s2726);
  and x930(s907,s1891,s511);
  and x931(s915,s1889,s505);
  and x932(s922,s1887,s499);
  and x933(s924,s493,s1885);
  and x934(s937,s1883,s540);
  and x935(s946,s1881,s534);
  or x936(s1109,s1107,s1108);
  and x937(s1125,s1953,s738);
  and x938(s1133,s1951,s732);
  and x939(s1140,s1949,s726);
  and x940(s1142,s720,s1947);
  and x941(s1155,s1945,s714);
  and x942(s1164,s1943,s708);
  or x943(s1378,s1368,s1369);
  or x944(s1380,s1371,s1373);
  or x945(s1382,s1375,s1377);
  or x946(s1624,s1614,s1615);
  or x947(s1626,s1617,s1619);
  or x948(s1628,s1621,s1623);
  not x949(s2725,s2719);
  or x950(s1859,s1856,s1858);
  or x951(s1864,s1861,s1863);
  or x952(s1921,s1918,s1920);
  or x953(s1926,s1923,s1925);
  buf x954(s2267,s1891);
  buf x955(s2275,s1889);
  buf x956(s2283,s1887);
  buf x957(s2291,s1885);
  buf x958(s2299,s1883);
  buf x959(s2307,s1881);
  buf x960(s2318,s528);
  buf x961(s2326,s522);
  buf x962(s2355,s1953);
  buf x963(s2363,s1951);
  buf x964(s2371,s1949);
  buf x965(s2379,s1947);
  buf x966(s2387,s1945);
  buf x967(s2395,s1943);
  buf x968(s2406,s702);
  buf x969(s2414,s696);
  nand x970(s647,s645,s646);
  nor x971(s631,s629,s630);
  nor x972(s634,s632,s633);
  nor x973(s637,s635,s636);
  nor x974(s640,s638,s639);
  not x975(s2234,s2230);
  not x976(s2250,s2246);
  and x977(s679,s677,s1031);
  nand x978(s1826,s2722,s2725);
  not x979(s2274,s2270);
  not x980(s2282,s2278);
  not x981(s2290,s2286);
  not x982(s2298,s2294);
  not x983(s2306,s2302);
  not x984(s2314,s2310);
  and x985(s1110,s1109,s1031);
  not x986(s2362,s2358);
  not x987(s2370,s2366);
  not x988(s2378,s2374);
  not x989(s2386,s2382);
  not x990(s2394,s2390);
  not x991(s2402,s2398);
  and x992(s1877,s1859,s1831);
  and x993(s1879,s1864,s1831);
  and x994(s1939,s1921,s1893);
  and x995(s1941,s1926,s1893);
  and x996(s143,s647,s865);
  and x997(s671,s1380,s1043);
  and x998(s674,s1378,s1035);
  nand x999(s686,s1826,s1827);
  not x1000(s2273,s2267);
  nand x1001(s900,s2267,s2274);
  not x1002(s2281,s2275);
  nand x1003(s909,s2275,s2282);
  not x1004(s2289,s2283);
  nand x1005(s917,s2283,s2290);
  not x1006(s2297,s2291);
  nand x1007(s926,s2291,s2298);
  not x1008(s2305,s2299);
  nand x1009(s929,s2299,s2306);
  not x1010(s2313,s2307);
  nand x1011(s939,s2307,s2314);
  not x1012(s2322,s2318);
  not x1013(s2330,s2326);
  and x1014(s967,s1382,s1051);
  and x1015(s1104,s1626,s1043);
  and x1016(s1106,s1624,s1035);
  not x1017(s2361,s2355);
  nand x1018(s1118,s2355,s2362);
  not x1019(s2369,s2363);
  nand x1020(s1127,s2363,s2370);
  not x1021(s2377,s2371);
  nand x1022(s1135,s2371,s2378);
  not x1023(s2385,s2379);
  nand x1024(s1144,s2379,s2386);
  not x1025(s2393,s2387);
  nand x1026(s1147,s2387,s2394);
  not x1027(s2401,s2395);
  nand x1028(s1157,s2395,s2402);
  not x1029(s2410,s2406);
  not x1030(s2418,s2414);
  and x1031(s1184,s1628,s1051);
  nand x1032(s2227,s634,s631);
  nand x1033(s2243,s640,s637);
  buf x1034(s2251,s1380);
  buf x1035(s2259,s1378);
  buf x1036(s2331,s1382);
  buf x1037(s2339,s1626);
  buf x1038(s2347,s1624);
  buf x1039(s2419,s1628);
  or x1040(s145,s143,s144);
  not x1041(s687,s686);
  nand x1042(s899,s2270,s2273);
  nand x1043(s908,s2278,s2281);
  nand x1044(s916,s2286,s2289);
  nand x1045(s925,s2294,s2297);
  nand x1046(s928,s2302,s2305);
  nand x1047(s938,s2310,s2313);
  and x1048(s954,s1879,s528);
  and x1049(s961,s1877,s522);
  nand x1050(s1117,s2358,s2361);
  nand x1051(s1126,s2366,s2369);
  nand x1052(s1134,s2374,s2377);
  nand x1053(s1143,s2382,s2385);
  nand x1054(s1146,s2390,s2393);
  nand x1055(s1156,s2398,s2401);
  and x1056(s1172,s1941,s702);
  and x1057(s1179,s1939,s696);
  buf x1058(s2315,s1879);
  buf x1059(s2323,s1877);
  buf x1060(s2403,s1941);
  buf x1061(s2411,s1939);
  not x1062(s2233,s2227);
  nand x1063(s642,s2227,s2234);
  not x1064(s2249,s2243);
  nand x1065(s649,s2243,s2250);
  not x1066(s2257,s2251);
  nand x1067(s665,s2251,s2258);
  nand x1068(s684,s2259,s2266);
  not x1069(s2265,s2259);
  and x1070(s688,s687,s487);
  nand x1071(s901,s899,s900);
  nand x1072(s910,s908,s909);
  nand x1073(s918,s916,s917);
  nand x1074(s927,s925,s926);
  nand x1075(s930,s928,s929);
  nand x1076(s940,s938,s939);
  not x1077(s2337,s2331);
  nand x1078(s963,s2331,s2338);
  not x1079(s2345,s2339);
  nand x1080(s1099,s2339,s2346);
  nand x1081(s1115,s2347,s2354);
  not x1082(s2353,s2347);
  nand x1083(s1119,s1117,s1118);
  nand x1084(s1128,s1126,s1127);
  nand x1085(s1136,s1134,s1135);
  nand x1086(s1145,s1143,s1144);
  nand x1087(s1148,s1146,s1147);
  nand x1088(s1158,s1156,s1157);
  not x1089(s2425,s2419);
  nand x1090(s1181,s2419,s2426);
  nand x1091(s641,s2230,s2233);
  nand x1092(s648,s2246,s2249);
  nand x1093(s664,s2254,s2257);
  nand x1094(s683,s2262,s2265);
  buf x1095(s395,s688);
  not x1096(s2321,s2315);
  nand x1097(s948,s2315,s2322);
  not x1098(s2329,s2323);
  nand x1099(s956,s2323,s2330);
  nand x1100(s962,s2334,s2337);
  nand x1101(s1098,s2342,s2345);
  nand x1102(s1114,s2350,s2353);
  not x1103(s2409,s2403);
  nand x1104(s1166,s2403,s2410);
  not x1105(s2417,s2411);
  nand x1106(s1174,s2411,s2418);
  nand x1107(s1180,s2422,s2425);
  nand x1108(s643,s641,s642);
  nand x1109(s650,s648,s649);
  nand x1110(s666,s664,s665);
  nand x1111(s681,s683,s684);
  not x1112(s690,s688);
  nand x1113(s947,s2318,s2321);
  nand x1114(s955,s2326,s2329);
  nand x1115(s964,s962,s963);
  and x1116(s968,s910,s927,s918,s901);
  and x1117(s970,s901,s915);
  and x1118(s971,s910,s901,s922);
  and x1119(s972,s918,s901,s924,s910);
  and x1120(s978,s930,s946);
  and x1121(s979,s940,s930,s954);
  nand x1122(s1100,s1098,s1099);
  nand x1123(s1112,s1114,s1115);
  nand x1124(s1165,s2406,s2409);
  nand x1125(s1173,s2414,s2417);
  nand x1126(s1182,s1180,s1181);
  and x1127(s1185,s1128,s1145,s1136,s1119);
  and x1128(s1187,s1119,s1133);
  and x1129(s1188,s1128,s1119,s1140);
  and x1130(s1189,s1136,s1119,s1142,s1128);
  and x1131(s1195,s1148,s1164);
  and x1132(s1196,s1158,s1148,s1172);
  not x1133(s644,s643);
  and x1134(s884,s650,s868);
  nand x1135(s949,s947,s948);
  nand x1136(s957,s955,s956);
  not x1137(s969,s968);
  or x1138(s973,s907,s970,s971,s972);
  nand x1139(s1167,s1165,s1166);
  nand x1140(s1175,s1173,s1174);
  not x1141(s1186,s1185);
  or x1142(s1190,s1125,s1187,s1188,s1189);
  and x1143(s680,s666,s674);
  and x1144(s682,s681,s666,s679);
  or x1145(s895,s883,s884);
  and x1146(s1025,s644,s487);
  and x1147(s1111,s1100,s1106);
  and x1148(s1113,s1112,s1100,s1110);
  or x1149(s685,s671,s680,s682);
  buf x1150(s295,s895);
  buf x1151(s331,s895);
  not x1152(s976,s973);
  and x1153(s977,s940,s964,s949,s930,s957);
  and x1154(s980,s949,s930,s961,s940);
  and x1155(s981,s957,s949,s930,s967,s940);
  buf x1156(s397,s1025);
  or x1157(s1116,s1104,s1111,s1113);
  not x1158(s1193,s1190);
  and x1159(s1194,s1158,s1182,s1167,s1148,s1175);
  and x1160(s1197,s1167,s1148,s1179,s1158);
  and x1161(s1198,s1175,s1167,s1148,s1184,s1158);
  or x1162(s982,s937,s978,s979,s980,s981);
  and x1163(s983,s977,s685);
  nand x1164(s988,s976,s969);
  not x1165(s1027,s1025);
  or x1166(s1199,s1155,s1195,s1196,s1197,s1198);
  and x1167(s1200,s1194,s1116);
  nand x1168(s1205,s1193,s1186);
  or x1169(s984,s982,s983);
  and x1170(s1085,s690,s1027,s1830);
  or x1171(s1201,s1199,s1200);
  not x1172(s987,s984);
  and x1173(s990,s988,s984);
  not x1174(s1204,s1201);
  and x1175(s1207,s1205,s1201);
  and x1176(s989,s973,s987);
  and x1177(s1206,s1190,s1204);
  or x1178(s991,s989,s990);
  or x1179(s1208,s1206,s1207);
  buf x1180(s329,s1208);
  nand x1181(s1221,s1208,s991);
  and x1182(s1238,s1208,s1221);
  and x1183(s1239,s1221,s991);
  or x1184(s1240,s1238,s1239);
  not x1185(s1247,s1240);
  and x1186(s471,s1240,s1247);
  or x1187(s473,s471,s1247);
  not x1188(s231,s473);
  and x1189(s1088,s1553,s1087,s473);
  and x1190(s1089,s1085,s1088,s554);
  buf x1191(s308,s1089);
  not x1192(s225,s1089);

endmodule
