module c1355(s1324gat,s1325gat,s1326gat,s1327gat,s1328gat,s1329gat,s1330gat,s1331gat,s1332gat,s1333gat,s1334gat,s1335gat,s1336gat,s1337gat,s1338gat,s1339gat,s1340gat,s1341gat,s1342gat,s1343gat,s1344gat,s1345gat,s1346gat,s1347gat,s1348gat,s1349gat,s1350gat,s1351gat,s1352gat,s1353gat,s1354gat,s1355gat,s1gat,s8gat,s15gat,s22gat,s29gat,s36gat,s43gat,s50gat,s57gat,s64gat,s71gat,s78gat,s85gat,s92gat,s99gat,s106gat,s113gat,s120gat,s127gat,s134gat,s141gat,s148gat,s155gat,s162gat,s169gat,s176gat,s183gat,s190gat,s197gat,s204gat,s211gat,s218gat,s225gat,s226gat,s227gat,s228gat,s229gat,s230gat,s231gat,s232gat,s233gat);

  output s1324gat;
  output s1325gat;
  output s1326gat;
  output s1327gat;
  output s1328gat;
  output s1329gat;
  output s1330gat;
  output s1331gat;
  output s1332gat;
  output s1333gat;
  output s1334gat;
  output s1335gat;
  output s1336gat;
  output s1337gat;
  output s1338gat;
  output s1339gat;
  output s1340gat;
  output s1341gat;
  output s1342gat;
  output s1343gat;
  output s1344gat;
  output s1345gat;
  output s1346gat;
  output s1347gat;
  output s1348gat;
  output s1349gat;
  output s1350gat;
  output s1351gat;
  output s1352gat;
  output s1353gat;
  output s1354gat;
  output s1355gat;
  input s1gat;
  input s8gat;
  input s15gat;
  input s22gat;
  input s29gat;
  input s36gat;
  input s43gat;
  input s50gat;
  input s57gat;
  input s64gat;
  input s71gat;
  input s78gat;
  input s85gat;
  input s92gat;
  input s99gat;
  input s106gat;
  input s113gat;
  input s120gat;
  input s127gat;
  input s134gat;
  input s141gat;
  input s148gat;
  input s155gat;
  input s162gat;
  input s169gat;
  input s176gat;
  input s183gat;
  input s190gat;
  input s197gat;
  input s204gat;
  input s211gat;
  input s218gat;
  input s225gat;
  input s226gat;
  input s227gat;
  input s228gat;
  input s229gat;
  input s230gat;
  input s231gat;
  input s232gat;
  input s233gat;

  and x0(s242gat,s225gat,s233gat);
  and x1(s245gat,s226gat,s233gat);
  and x2(s248gat,s227gat,s233gat);
  and x3(s251gat,s228gat,s233gat);
  and x4(s254gat,s229gat,s233gat);
  and x5(s257gat,s230gat,s233gat);
  and x6(s260gat,s231gat,s233gat);
  and x7(s263gat,s232gat,s233gat);
  nand x8(s266gat,s1gat,s8gat);
  nand x9(s269gat,s15gat,s22gat);
  nand x10(s272gat,s29gat,s36gat);
  nand x11(s275gat,s43gat,s50gat);
  nand x12(s278gat,s57gat,s64gat);
  nand x13(s281gat,s71gat,s78gat);
  nand x14(s284gat,s85gat,s92gat);
  nand x15(s287gat,s99gat,s106gat);
  nand x16(s290gat,s113gat,s120gat);
  nand x17(s293gat,s127gat,s134gat);
  nand x18(s296gat,s141gat,s148gat);
  nand x19(s299gat,s155gat,s162gat);
  nand x20(s302gat,s169gat,s176gat);
  nand x21(s305gat,s183gat,s190gat);
  nand x22(s308gat,s197gat,s204gat);
  nand x23(s311gat,s211gat,s218gat);
  nand x24(s314gat,s1gat,s29gat);
  nand x25(s317gat,s57gat,s85gat);
  nand x26(s320gat,s8gat,s36gat);
  nand x27(s323gat,s64gat,s92gat);
  nand x28(s326gat,s15gat,s43gat);
  nand x29(s329gat,s71gat,s99gat);
  nand x30(s332gat,s22gat,s50gat);
  nand x31(s335gat,s78gat,s106gat);
  nand x32(s338gat,s113gat,s141gat);
  nand x33(s341gat,s169gat,s197gat);
  nand x34(s344gat,s120gat,s148gat);
  nand x35(s347gat,s176gat,s204gat);
  nand x36(s350gat,s127gat,s155gat);
  nand x37(s353gat,s183gat,s211gat);
  nand x38(s356gat,s134gat,s162gat);
  nand x39(s359gat,s190gat,s218gat);
  nand x40(s362gat,s1gat,s266gat);
  nand x41(s363gat,s8gat,s266gat);
  nand x42(s364gat,s15gat,s269gat);
  nand x43(s365gat,s22gat,s269gat);
  nand x44(s366gat,s29gat,s272gat);
  nand x45(s367gat,s36gat,s272gat);
  nand x46(s368gat,s43gat,s275gat);
  nand x47(s369gat,s50gat,s275gat);
  nand x48(s370gat,s57gat,s278gat);
  nand x49(s371gat,s64gat,s278gat);
  nand x50(s372gat,s71gat,s281gat);
  nand x51(s373gat,s78gat,s281gat);
  nand x52(s374gat,s85gat,s284gat);
  nand x53(s375gat,s92gat,s284gat);
  nand x54(s376gat,s99gat,s287gat);
  nand x55(s377gat,s106gat,s287gat);
  nand x56(s378gat,s113gat,s290gat);
  nand x57(s379gat,s120gat,s290gat);
  nand x58(s380gat,s127gat,s293gat);
  nand x59(s381gat,s134gat,s293gat);
  nand x60(s382gat,s141gat,s296gat);
  nand x61(s383gat,s148gat,s296gat);
  nand x62(s384gat,s155gat,s299gat);
  nand x63(s385gat,s162gat,s299gat);
  nand x64(s386gat,s169gat,s302gat);
  nand x65(s387gat,s176gat,s302gat);
  nand x66(s388gat,s183gat,s305gat);
  nand x67(s389gat,s190gat,s305gat);
  nand x68(s390gat,s197gat,s308gat);
  nand x69(s391gat,s204gat,s308gat);
  nand x70(s392gat,s211gat,s311gat);
  nand x71(s393gat,s218gat,s311gat);
  nand x72(s394gat,s1gat,s314gat);
  nand x73(s395gat,s29gat,s314gat);
  nand x74(s396gat,s57gat,s317gat);
  nand x75(s397gat,s85gat,s317gat);
  nand x76(s398gat,s8gat,s320gat);
  nand x77(s399gat,s36gat,s320gat);
  nand x78(s400gat,s64gat,s323gat);
  nand x79(s401gat,s92gat,s323gat);
  nand x80(s402gat,s15gat,s326gat);
  nand x81(s403gat,s43gat,s326gat);
  nand x82(s404gat,s71gat,s329gat);
  nand x83(s405gat,s99gat,s329gat);
  nand x84(s406gat,s22gat,s332gat);
  nand x85(s407gat,s50gat,s332gat);
  nand x86(s408gat,s78gat,s335gat);
  nand x87(s409gat,s106gat,s335gat);
  nand x88(s410gat,s113gat,s338gat);
  nand x89(s411gat,s141gat,s338gat);
  nand x90(s412gat,s169gat,s341gat);
  nand x91(s413gat,s197gat,s341gat);
  nand x92(s414gat,s120gat,s344gat);
  nand x93(s415gat,s148gat,s344gat);
  nand x94(s416gat,s176gat,s347gat);
  nand x95(s417gat,s204gat,s347gat);
  nand x96(s418gat,s127gat,s350gat);
  nand x97(s419gat,s155gat,s350gat);
  nand x98(s420gat,s183gat,s353gat);
  nand x99(s421gat,s211gat,s353gat);
  nand x100(s422gat,s134gat,s356gat);
  nand x101(s423gat,s162gat,s356gat);
  nand x102(s424gat,s190gat,s359gat);
  nand x103(s425gat,s218gat,s359gat);
  nand x104(s426gat,s362gat,s363gat);
  nand x105(s429gat,s364gat,s365gat);
  nand x106(s432gat,s366gat,s367gat);
  nand x107(s435gat,s368gat,s369gat);
  nand x108(s438gat,s370gat,s371gat);
  nand x109(s441gat,s372gat,s373gat);
  nand x110(s444gat,s374gat,s375gat);
  nand x111(s447gat,s376gat,s377gat);
  nand x112(s450gat,s378gat,s379gat);
  nand x113(s453gat,s380gat,s381gat);
  nand x114(s456gat,s382gat,s383gat);
  nand x115(s459gat,s384gat,s385gat);
  nand x116(s462gat,s386gat,s387gat);
  nand x117(s465gat,s388gat,s389gat);
  nand x118(s468gat,s390gat,s391gat);
  nand x119(s471gat,s392gat,s393gat);
  nand x120(s474gat,s394gat,s395gat);
  nand x121(s477gat,s396gat,s397gat);
  nand x122(s480gat,s398gat,s399gat);
  nand x123(s483gat,s400gat,s401gat);
  nand x124(s486gat,s402gat,s403gat);
  nand x125(s489gat,s404gat,s405gat);
  nand x126(s492gat,s406gat,s407gat);
  nand x127(s495gat,s408gat,s409gat);
  nand x128(s498gat,s410gat,s411gat);
  nand x129(s501gat,s412gat,s413gat);
  nand x130(s504gat,s414gat,s415gat);
  nand x131(s507gat,s416gat,s417gat);
  nand x132(s510gat,s418gat,s419gat);
  nand x133(s513gat,s420gat,s421gat);
  nand x134(s516gat,s422gat,s423gat);
  nand x135(s519gat,s424gat,s425gat);
  nand x136(s522gat,s426gat,s429gat);
  nand x137(s525gat,s432gat,s435gat);
  nand x138(s528gat,s438gat,s441gat);
  nand x139(s531gat,s444gat,s447gat);
  nand x140(s534gat,s450gat,s453gat);
  nand x141(s537gat,s456gat,s459gat);
  nand x142(s540gat,s462gat,s465gat);
  nand x143(s543gat,s468gat,s471gat);
  nand x144(s546gat,s474gat,s477gat);
  nand x145(s549gat,s480gat,s483gat);
  nand x146(s552gat,s486gat,s489gat);
  nand x147(s555gat,s492gat,s495gat);
  nand x148(s558gat,s498gat,s501gat);
  nand x149(s561gat,s504gat,s507gat);
  nand x150(s564gat,s510gat,s513gat);
  nand x151(s567gat,s516gat,s519gat);
  nand x152(s570gat,s426gat,s522gat);
  nand x153(s571gat,s429gat,s522gat);
  nand x154(s572gat,s432gat,s525gat);
  nand x155(s573gat,s435gat,s525gat);
  nand x156(s574gat,s438gat,s528gat);
  nand x157(s575gat,s441gat,s528gat);
  nand x158(s576gat,s444gat,s531gat);
  nand x159(s577gat,s447gat,s531gat);
  nand x160(s578gat,s450gat,s534gat);
  nand x161(s579gat,s453gat,s534gat);
  nand x162(s580gat,s456gat,s537gat);
  nand x163(s581gat,s459gat,s537gat);
  nand x164(s582gat,s462gat,s540gat);
  nand x165(s583gat,s465gat,s540gat);
  nand x166(s584gat,s468gat,s543gat);
  nand x167(s585gat,s471gat,s543gat);
  nand x168(s586gat,s474gat,s546gat);
  nand x169(s587gat,s477gat,s546gat);
  nand x170(s588gat,s480gat,s549gat);
  nand x171(s589gat,s483gat,s549gat);
  nand x172(s590gat,s486gat,s552gat);
  nand x173(s591gat,s489gat,s552gat);
  nand x174(s592gat,s492gat,s555gat);
  nand x175(s593gat,s495gat,s555gat);
  nand x176(s594gat,s498gat,s558gat);
  nand x177(s595gat,s501gat,s558gat);
  nand x178(s596gat,s504gat,s561gat);
  nand x179(s597gat,s507gat,s561gat);
  nand x180(s598gat,s510gat,s564gat);
  nand x181(s599gat,s513gat,s564gat);
  nand x182(s600gat,s516gat,s567gat);
  nand x183(s601gat,s519gat,s567gat);
  nand x184(s602gat,s570gat,s571gat);
  nand x185(s607gat,s572gat,s573gat);
  nand x186(s612gat,s574gat,s575gat);
  nand x187(s617gat,s576gat,s577gat);
  nand x188(s622gat,s578gat,s579gat);
  nand x189(s627gat,s580gat,s581gat);
  nand x190(s632gat,s582gat,s583gat);
  nand x191(s637gat,s584gat,s585gat);
  nand x192(s642gat,s586gat,s587gat);
  nand x193(s645gat,s588gat,s589gat);
  nand x194(s648gat,s590gat,s591gat);
  nand x195(s651gat,s592gat,s593gat);
  nand x196(s654gat,s594gat,s595gat);
  nand x197(s657gat,s596gat,s597gat);
  nand x198(s660gat,s598gat,s599gat);
  nand x199(s663gat,s600gat,s601gat);
  nand x200(s666gat,s602gat,s607gat);
  nand x201(s669gat,s612gat,s617gat);
  nand x202(s672gat,s602gat,s612gat);
  nand x203(s675gat,s607gat,s617gat);
  nand x204(s678gat,s622gat,s627gat);
  nand x205(s681gat,s632gat,s637gat);
  nand x206(s684gat,s622gat,s632gat);
  nand x207(s687gat,s627gat,s637gat);
  nand x208(s690gat,s602gat,s666gat);
  nand x209(s691gat,s607gat,s666gat);
  nand x210(s692gat,s612gat,s669gat);
  nand x211(s693gat,s617gat,s669gat);
  nand x212(s694gat,s602gat,s672gat);
  nand x213(s695gat,s612gat,s672gat);
  nand x214(s696gat,s607gat,s675gat);
  nand x215(s697gat,s617gat,s675gat);
  nand x216(s698gat,s622gat,s678gat);
  nand x217(s699gat,s627gat,s678gat);
  nand x218(s700gat,s632gat,s681gat);
  nand x219(s701gat,s637gat,s681gat);
  nand x220(s702gat,s622gat,s684gat);
  nand x221(s703gat,s632gat,s684gat);
  nand x222(s704gat,s627gat,s687gat);
  nand x223(s705gat,s637gat,s687gat);
  nand x224(s706gat,s690gat,s691gat);
  nand x225(s709gat,s692gat,s693gat);
  nand x226(s712gat,s694gat,s695gat);
  nand x227(s715gat,s696gat,s697gat);
  nand x228(s718gat,s698gat,s699gat);
  nand x229(s721gat,s700gat,s701gat);
  nand x230(s724gat,s702gat,s703gat);
  nand x231(s727gat,s704gat,s705gat);
  nand x232(s730gat,s242gat,s718gat);
  nand x233(s733gat,s245gat,s721gat);
  nand x234(s736gat,s248gat,s724gat);
  nand x235(s739gat,s251gat,s727gat);
  nand x236(s742gat,s254gat,s706gat);
  nand x237(s745gat,s257gat,s709gat);
  nand x238(s748gat,s260gat,s712gat);
  nand x239(s751gat,s263gat,s715gat);
  nand x240(s754gat,s242gat,s730gat);
  nand x241(s755gat,s718gat,s730gat);
  nand x242(s756gat,s245gat,s733gat);
  nand x243(s757gat,s721gat,s733gat);
  nand x244(s758gat,s248gat,s736gat);
  nand x245(s759gat,s724gat,s736gat);
  nand x246(s760gat,s251gat,s739gat);
  nand x247(s761gat,s727gat,s739gat);
  nand x248(s762gat,s254gat,s742gat);
  nand x249(s763gat,s706gat,s742gat);
  nand x250(s764gat,s257gat,s745gat);
  nand x251(s765gat,s709gat,s745gat);
  nand x252(s766gat,s260gat,s748gat);
  nand x253(s767gat,s712gat,s748gat);
  nand x254(s768gat,s263gat,s751gat);
  nand x255(s769gat,s715gat,s751gat);
  nand x256(s770gat,s754gat,s755gat);
  nand x257(s773gat,s756gat,s757gat);
  nand x258(s776gat,s758gat,s759gat);
  nand x259(s779gat,s760gat,s761gat);
  nand x260(s782gat,s762gat,s763gat);
  nand x261(s785gat,s764gat,s765gat);
  nand x262(s788gat,s766gat,s767gat);
  nand x263(s791gat,s768gat,s769gat);
  nand x264(s794gat,s642gat,s770gat);
  nand x265(s797gat,s645gat,s773gat);
  nand x266(s800gat,s648gat,s776gat);
  nand x267(s803gat,s651gat,s779gat);
  nand x268(s806gat,s654gat,s782gat);
  nand x269(s809gat,s657gat,s785gat);
  nand x270(s812gat,s660gat,s788gat);
  nand x271(s815gat,s663gat,s791gat);
  nand x272(s818gat,s642gat,s794gat);
  nand x273(s819gat,s770gat,s794gat);
  nand x274(s820gat,s645gat,s797gat);
  nand x275(s821gat,s773gat,s797gat);
  nand x276(s822gat,s648gat,s800gat);
  nand x277(s823gat,s776gat,s800gat);
  nand x278(s824gat,s651gat,s803gat);
  nand x279(s825gat,s779gat,s803gat);
  nand x280(s826gat,s654gat,s806gat);
  nand x281(s827gat,s782gat,s806gat);
  nand x282(s828gat,s657gat,s809gat);
  nand x283(s829gat,s785gat,s809gat);
  nand x284(s830gat,s660gat,s812gat);
  nand x285(s831gat,s788gat,s812gat);
  nand x286(s832gat,s663gat,s815gat);
  nand x287(s833gat,s791gat,s815gat);
  nand x288(s834gat,s818gat,s819gat);
  nand x289(s847gat,s820gat,s821gat);
  nand x290(s860gat,s822gat,s823gat);
  nand x291(s873gat,s824gat,s825gat);
  nand x292(s886gat,s828gat,s829gat);
  nand x293(s899gat,s832gat,s833gat);
  nand x294(s912gat,s830gat,s831gat);
  nand x295(s925gat,s826gat,s827gat);
  not x296(s938gat,s834gat);
  not x297(s939gat,s847gat);
  not x298(s940gat,s860gat);
  not x299(s941gat,s834gat);
  not x300(s942gat,s847gat);
  not x301(s943gat,s873gat);
  not x302(s944gat,s834gat);
  not x303(s945gat,s860gat);
  not x304(s946gat,s873gat);
  not x305(s947gat,s847gat);
  not x306(s948gat,s860gat);
  not x307(s949gat,s873gat);
  not x308(s950gat,s886gat);
  not x309(s951gat,s899gat);
  not x310(s952gat,s886gat);
  not x311(s953gat,s912gat);
  not x312(s954gat,s925gat);
  not x313(s955gat,s899gat);
  not x314(s956gat,s925gat);
  not x315(s957gat,s912gat);
  not x316(s958gat,s925gat);
  not x317(s959gat,s886gat);
  not x318(s960gat,s912gat);
  not x319(s961gat,s925gat);
  not x320(s962gat,s886gat);
  not x321(s963gat,s899gat);
  not x322(s964gat,s925gat);
  not x323(s965gat,s912gat);
  not x324(s966gat,s899gat);
  not x325(s967gat,s886gat);
  not x326(s968gat,s912gat);
  not x327(s969gat,s899gat);
  not x328(s970gat,s847gat);
  not x329(s971gat,s873gat);
  not x330(s972gat,s847gat);
  not x331(s973gat,s860gat);
  not x332(s974gat,s834gat);
  not x333(s975gat,s873gat);
  not x334(s976gat,s834gat);
  not x335(s977gat,s860gat);
  and x336(s978gat,s938gat,s939gat,s940gat,s873gat);
  and x337(s979gat,s941gat,s942gat,s860gat,s943gat);
  and x338(s980gat,s944gat,s847gat,s945gat,s946gat);
  and x339(s981gat,s834gat,s947gat,s948gat,s949gat);
  and x340(s982gat,s958gat,s959gat,s960gat,s899gat);
  and x341(s983gat,s961gat,s962gat,s912gat,s963gat);
  and x342(s984gat,s964gat,s886gat,s965gat,s966gat);
  and x343(s985gat,s925gat,s967gat,s968gat,s969gat);
  or x344(s986gat,s978gat,s979gat,s980gat,s981gat);
  or x345(s991gat,s982gat,s983gat,s984gat,s985gat);
  and x346(s996gat,s925gat,s950gat,s912gat,s951gat,s986gat);
  and x347(s1001gat,s925gat,s952gat,s953gat,s899gat,s986gat);
  and x348(s1006gat,s954gat,s886gat,s912gat,s955gat,s986gat);
  and x349(s1011gat,s956gat,s886gat,s957gat,s899gat,s986gat);
  and x350(s1016gat,s834gat,s970gat,s860gat,s971gat,s991gat);
  and x351(s1021gat,s834gat,s972gat,s973gat,s873gat,s991gat);
  and x352(s1026gat,s974gat,s847gat,s860gat,s975gat,s991gat);
  and x353(s1031gat,s976gat,s847gat,s977gat,s873gat,s991gat);
  and x354(s1036gat,s834gat,s996gat);
  and x355(s1039gat,s847gat,s996gat);
  and x356(s1042gat,s860gat,s996gat);
  and x357(s1045gat,s873gat,s996gat);
  and x358(s1048gat,s834gat,s1001gat);
  and x359(s1051gat,s847gat,s1001gat);
  and x360(s1054gat,s860gat,s1001gat);
  and x361(s1057gat,s873gat,s1001gat);
  and x362(s1060gat,s834gat,s1006gat);
  and x363(s1063gat,s847gat,s1006gat);
  and x364(s1066gat,s860gat,s1006gat);
  and x365(s1069gat,s873gat,s1006gat);
  and x366(s1072gat,s834gat,s1011gat);
  and x367(s1075gat,s847gat,s1011gat);
  and x368(s1078gat,s860gat,s1011gat);
  and x369(s1081gat,s873gat,s1011gat);
  and x370(s1084gat,s925gat,s1016gat);
  and x371(s1087gat,s886gat,s1016gat);
  and x372(s1090gat,s912gat,s1016gat);
  and x373(s1093gat,s899gat,s1016gat);
  and x374(s1096gat,s925gat,s1021gat);
  and x375(s1099gat,s886gat,s1021gat);
  and x376(s1102gat,s912gat,s1021gat);
  and x377(s1105gat,s899gat,s1021gat);
  and x378(s1108gat,s925gat,s1026gat);
  and x379(s1111gat,s886gat,s1026gat);
  and x380(s1114gat,s912gat,s1026gat);
  and x381(s1117gat,s899gat,s1026gat);
  and x382(s1120gat,s925gat,s1031gat);
  and x383(s1123gat,s886gat,s1031gat);
  and x384(s1126gat,s912gat,s1031gat);
  and x385(s1129gat,s899gat,s1031gat);
  nand x386(s1132gat,s1gat,s1036gat);
  nand x387(s1135gat,s8gat,s1039gat);
  nand x388(s1138gat,s15gat,s1042gat);
  nand x389(s1141gat,s22gat,s1045gat);
  nand x390(s1144gat,s29gat,s1048gat);
  nand x391(s1147gat,s36gat,s1051gat);
  nand x392(s1150gat,s43gat,s1054gat);
  nand x393(s1153gat,s50gat,s1057gat);
  nand x394(s1156gat,s57gat,s1060gat);
  nand x395(s1159gat,s64gat,s1063gat);
  nand x396(s1162gat,s71gat,s1066gat);
  nand x397(s1165gat,s78gat,s1069gat);
  nand x398(s1168gat,s85gat,s1072gat);
  nand x399(s1171gat,s92gat,s1075gat);
  nand x400(s1174gat,s99gat,s1078gat);
  nand x401(s1177gat,s106gat,s1081gat);
  nand x402(s1180gat,s113gat,s1084gat);
  nand x403(s1183gat,s120gat,s1087gat);
  nand x404(s1186gat,s127gat,s1090gat);
  nand x405(s1189gat,s134gat,s1093gat);
  nand x406(s1192gat,s141gat,s1096gat);
  nand x407(s1195gat,s148gat,s1099gat);
  nand x408(s1198gat,s155gat,s1102gat);
  nand x409(s1201gat,s162gat,s1105gat);
  nand x410(s1204gat,s169gat,s1108gat);
  nand x411(s1207gat,s176gat,s1111gat);
  nand x412(s1210gat,s183gat,s1114gat);
  nand x413(s1213gat,s190gat,s1117gat);
  nand x414(s1216gat,s197gat,s1120gat);
  nand x415(s1219gat,s204gat,s1123gat);
  nand x416(s1222gat,s211gat,s1126gat);
  nand x417(s1225gat,s218gat,s1129gat);
  nand x418(s1228gat,s1gat,s1132gat);
  nand x419(s1229gat,s1036gat,s1132gat);
  nand x420(s1230gat,s8gat,s1135gat);
  nand x421(s1231gat,s1039gat,s1135gat);
  nand x422(s1232gat,s15gat,s1138gat);
  nand x423(s1233gat,s1042gat,s1138gat);
  nand x424(s1234gat,s22gat,s1141gat);
  nand x425(s1235gat,s1045gat,s1141gat);
  nand x426(s1236gat,s29gat,s1144gat);
  nand x427(s1237gat,s1048gat,s1144gat);
  nand x428(s1238gat,s36gat,s1147gat);
  nand x429(s1239gat,s1051gat,s1147gat);
  nand x430(s1240gat,s43gat,s1150gat);
  nand x431(s1241gat,s1054gat,s1150gat);
  nand x432(s1242gat,s50gat,s1153gat);
  nand x433(s1243gat,s1057gat,s1153gat);
  nand x434(s1244gat,s57gat,s1156gat);
  nand x435(s1245gat,s1060gat,s1156gat);
  nand x436(s1246gat,s64gat,s1159gat);
  nand x437(s1247gat,s1063gat,s1159gat);
  nand x438(s1248gat,s71gat,s1162gat);
  nand x439(s1249gat,s1066gat,s1162gat);
  nand x440(s1250gat,s78gat,s1165gat);
  nand x441(s1251gat,s1069gat,s1165gat);
  nand x442(s1252gat,s85gat,s1168gat);
  nand x443(s1253gat,s1072gat,s1168gat);
  nand x444(s1254gat,s92gat,s1171gat);
  nand x445(s1255gat,s1075gat,s1171gat);
  nand x446(s1256gat,s99gat,s1174gat);
  nand x447(s1257gat,s1078gat,s1174gat);
  nand x448(s1258gat,s106gat,s1177gat);
  nand x449(s1259gat,s1081gat,s1177gat);
  nand x450(s1260gat,s113gat,s1180gat);
  nand x451(s1261gat,s1084gat,s1180gat);
  nand x452(s1262gat,s120gat,s1183gat);
  nand x453(s1263gat,s1087gat,s1183gat);
  nand x454(s1264gat,s127gat,s1186gat);
  nand x455(s1265gat,s1090gat,s1186gat);
  nand x456(s1266gat,s134gat,s1189gat);
  nand x457(s1267gat,s1093gat,s1189gat);
  nand x458(s1268gat,s141gat,s1192gat);
  nand x459(s1269gat,s1096gat,s1192gat);
  nand x460(s1270gat,s148gat,s1195gat);
  nand x461(s1271gat,s1099gat,s1195gat);
  nand x462(s1272gat,s155gat,s1198gat);
  nand x463(s1273gat,s1102gat,s1198gat);
  nand x464(s1274gat,s162gat,s1201gat);
  nand x465(s1275gat,s1105gat,s1201gat);
  nand x466(s1276gat,s169gat,s1204gat);
  nand x467(s1277gat,s1108gat,s1204gat);
  nand x468(s1278gat,s176gat,s1207gat);
  nand x469(s1279gat,s1111gat,s1207gat);
  nand x470(s1280gat,s183gat,s1210gat);
  nand x471(s1281gat,s1114gat,s1210gat);
  nand x472(s1282gat,s190gat,s1213gat);
  nand x473(s1283gat,s1117gat,s1213gat);
  nand x474(s1284gat,s197gat,s1216gat);
  nand x475(s1285gat,s1120gat,s1216gat);
  nand x476(s1286gat,s204gat,s1219gat);
  nand x477(s1287gat,s1123gat,s1219gat);
  nand x478(s1288gat,s211gat,s1222gat);
  nand x479(s1289gat,s1126gat,s1222gat);
  nand x480(s1290gat,s218gat,s1225gat);
  nand x481(s1291gat,s1129gat,s1225gat);
  nand x482(s1292gat,s1228gat,s1229gat);
  nand x483(s1293gat,s1230gat,s1231gat);
  nand x484(s1294gat,s1232gat,s1233gat);
  nand x485(s1295gat,s1234gat,s1235gat);
  nand x486(s1296gat,s1236gat,s1237gat);
  nand x487(s1297gat,s1238gat,s1239gat);
  nand x488(s1298gat,s1240gat,s1241gat);
  nand x489(s1299gat,s1242gat,s1243gat);
  nand x490(s1300gat,s1244gat,s1245gat);
  nand x491(s1301gat,s1246gat,s1247gat);
  nand x492(s1302gat,s1248gat,s1249gat);
  nand x493(s1303gat,s1250gat,s1251gat);
  nand x494(s1304gat,s1252gat,s1253gat);
  nand x495(s1305gat,s1254gat,s1255gat);
  nand x496(s1306gat,s1256gat,s1257gat);
  nand x497(s1307gat,s1258gat,s1259gat);
  nand x498(s1308gat,s1260gat,s1261gat);
  nand x499(s1309gat,s1262gat,s1263gat);
  nand x500(s1310gat,s1264gat,s1265gat);
  nand x501(s1311gat,s1266gat,s1267gat);
  nand x502(s1312gat,s1268gat,s1269gat);
  nand x503(s1313gat,s1270gat,s1271gat);
  nand x504(s1314gat,s1272gat,s1273gat);
  nand x505(s1315gat,s1274gat,s1275gat);
  nand x506(s1316gat,s1276gat,s1277gat);
  nand x507(s1317gat,s1278gat,s1279gat);
  nand x508(s1318gat,s1280gat,s1281gat);
  nand x509(s1319gat,s1282gat,s1283gat);
  nand x510(s1320gat,s1284gat,s1285gat);
  nand x511(s1321gat,s1286gat,s1287gat);
  nand x512(s1322gat,s1288gat,s1289gat);
  nand x513(s1323gat,s1290gat,s1291gat);
  buf x514(s1324gat,s1292gat);
  buf x515(s1325gat,s1293gat);
  buf x516(s1326gat,s1294gat);
  buf x517(s1327gat,s1295gat);
  buf x518(s1328gat,s1296gat);
  buf x519(s1329gat,s1297gat);
  buf x520(s1330gat,s1298gat);
  buf x521(s1331gat,s1299gat);
  buf x522(s1332gat,s1300gat);
  buf x523(s1333gat,s1301gat);
  buf x524(s1334gat,s1302gat);
  buf x525(s1335gat,s1303gat);
  buf x526(s1336gat,s1304gat);
  buf x527(s1337gat,s1305gat);
  buf x528(s1338gat,s1306gat);
  buf x529(s1339gat,s1307gat);
  buf x530(s1340gat,s1308gat);
  buf x531(s1341gat,s1309gat);
  buf x532(s1342gat,s1310gat);
  buf x533(s1343gat,s1311gat);
  buf x534(s1344gat,s1312gat);
  buf x535(s1345gat,s1313gat);
  buf x536(s1346gat,s1314gat);
  buf x537(s1347gat,s1315gat);
  buf x538(s1348gat,s1316gat);
  buf x539(s1349gat,s1317gat);
  buf x540(s1350gat,s1318gat);
  buf x541(s1351gat,s1319gat);
  buf x542(s1352gat,s1320gat);
  buf x543(s1353gat,s1321gat);
  buf x544(s1354gat,s1322gat);
  buf x545(s1355gat,s1323gat);

endmodule
