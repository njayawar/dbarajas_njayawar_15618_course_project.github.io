module c880(s388gat,s389gat,s390gat,s391gat,s418gat,s419gat,s420gat,s421gat,s422gat,s423gat,s446gat,s447gat,s448gat,s449gat,s450gat,s767gat,s768gat,s850gat,s863gat,s864gat,s865gat,s866gat,s874gat,s878gat,s879gat,s880gat,s1gat,s8gat,s13gat,s17gat,s26gat,s29gat,s36gat,s42gat,s51gat,s55gat,s59gat,s68gat,s72gat,s73gat,s74gat,s75gat,s80gat,s85gat,s86gat,s87gat,s88gat,s89gat,s90gat,s91gat,s96gat,s101gat,s106gat,s111gat,s116gat,s121gat,s126gat,s130gat,s135gat,s138gat,s143gat,s146gat,s149gat,s152gat,s153gat,s156gat,s159gat,s165gat,s171gat,s177gat,s183gat,s189gat,s195gat,s201gat,s207gat,s210gat,s219gat,s228gat,s237gat,s246gat,s255gat,s259gat,s260gat,s261gat,s267gat,s268gat);

  output s388gat;
  output s389gat;
  output s390gat;
  output s391gat;
  output s418gat;
  output s419gat;
  output s420gat;
  output s421gat;
  output s422gat;
  output s423gat;
  output s446gat;
  output s447gat;
  output s448gat;
  output s449gat;
  output s450gat;
  output s767gat;
  output s768gat;
  output s850gat;
  output s863gat;
  output s864gat;
  output s865gat;
  output s866gat;
  output s874gat;
  output s878gat;
  output s879gat;
  output s880gat;
  input s1gat;
  input s8gat;
  input s13gat;
  input s17gat;
  input s26gat;
  input s29gat;
  input s36gat;
  input s42gat;
  input s51gat;
  input s55gat;
  input s59gat;
  input s68gat;
  input s72gat;
  input s73gat;
  input s74gat;
  input s75gat;
  input s80gat;
  input s85gat;
  input s86gat;
  input s87gat;
  input s88gat;
  input s89gat;
  input s90gat;
  input s91gat;
  input s96gat;
  input s101gat;
  input s106gat;
  input s111gat;
  input s116gat;
  input s121gat;
  input s126gat;
  input s130gat;
  input s135gat;
  input s138gat;
  input s143gat;
  input s146gat;
  input s149gat;
  input s152gat;
  input s153gat;
  input s156gat;
  input s159gat;
  input s165gat;
  input s171gat;
  input s177gat;
  input s183gat;
  input s189gat;
  input s195gat;
  input s201gat;
  input s207gat;
  input s210gat;
  input s219gat;
  input s228gat;
  input s237gat;
  input s246gat;
  input s255gat;
  input s259gat;
  input s260gat;
  input s261gat;
  input s267gat;
  input s268gat;

  nand x0(s269gat,s1gat,s8gat,s13gat,s17gat);
  nand x1(s270gat,s1gat,s26gat,s13gat,s17gat);
  and x2(s273gat,s29gat,s36gat,s42gat);
  and x3(s276gat,s1gat,s26gat,s51gat);
  nand x4(s279gat,s1gat,s8gat,s51gat,s17gat);
  nand x5(s280gat,s1gat,s8gat,s13gat,s55gat);
  nand x6(s284gat,s59gat,s42gat,s68gat,s72gat);
  nand x7(s285gat,s29gat,s68gat);
  nand x8(s286gat,s59gat,s68gat,s74gat);
  and x9(s287gat,s29gat,s75gat,s80gat);
  and x10(s290gat,s29gat,s75gat,s42gat);
  and x11(s291gat,s29gat,s36gat,s80gat);
  and x12(s292gat,s29gat,s36gat,s42gat);
  and x13(s293gat,s59gat,s75gat,s80gat);
  and x14(s294gat,s59gat,s75gat,s42gat);
  and x15(s295gat,s59gat,s36gat,s80gat);
  and x16(s296gat,s59gat,s36gat,s42gat);
  and x17(s297gat,s85gat,s86gat);
  or x18(s298gat,s87gat,s88gat);
  nand x19(s301gat,s91gat,s96gat);
  or x20(s302gat,s91gat,s96gat);
  nand x21(s303gat,s101gat,s106gat);
  or x22(s304gat,s101gat,s106gat);
  nand x23(s305gat,s111gat,s116gat);
  or x24(s306gat,s111gat,s116gat);
  nand x25(s307gat,s121gat,s126gat);
  or x26(s308gat,s121gat,s126gat);
  and x27(s309gat,s8gat,s138gat);
  not x28(s310gat,s268gat);
  and x29(s316gat,s51gat,s138gat);
  and x30(s317gat,s17gat,s138gat);
  and x31(s318gat,s152gat,s138gat);
  nand x32(s319gat,s59gat,s156gat);
  nor x33(s322gat,s17gat,s42gat);
  and x34(s323gat,s17gat,s42gat);
  nand x35(s324gat,s159gat,s165gat);
  or x36(s325gat,s159gat,s165gat);
  nand x37(s326gat,s171gat,s177gat);
  or x38(s327gat,s171gat,s177gat);
  nand x39(s328gat,s183gat,s189gat);
  or x40(s329gat,s183gat,s189gat);
  nand x41(s330gat,s195gat,s201gat);
  or x42(s331gat,s195gat,s201gat);
  and x43(s332gat,s210gat,s91gat);
  and x44(s333gat,s210gat,s96gat);
  and x45(s334gat,s210gat,s101gat);
  and x46(s335gat,s210gat,s106gat);
  and x47(s336gat,s210gat,s111gat);
  and x48(s337gat,s255gat,s259gat);
  and x49(s338gat,s210gat,s116gat);
  and x50(s339gat,s255gat,s260gat);
  and x51(s340gat,s210gat,s121gat);
  and x52(s341gat,s255gat,s267gat);
  not x53(s342gat,s269gat);
  not x54(s343gat,s273gat);
  or x55(s344gat,s270gat,s273gat);
  not x56(s345gat,s276gat);
  not x57(s346gat,s276gat);
  not x58(s347gat,s279gat);
  nor x59(s348gat,s280gat,s284gat);
  or x60(s349gat,s280gat,s285gat);
  or x61(s350gat,s280gat,s286gat);
  not x62(s351gat,s293gat);
  not x63(s352gat,s294gat);
  not x64(s353gat,s295gat);
  not x65(s354gat,s296gat);
  nand x66(s355gat,s89gat,s298gat);
  and x67(s356gat,s90gat,s298gat);
  nand x68(s357gat,s301gat,s302gat);
  nand x69(s360gat,s303gat,s304gat);
  nand x70(s363gat,s305gat,s306gat);
  nand x71(s366gat,s307gat,s308gat);
  not x72(s369gat,s310gat);
  nor x73(s375gat,s322gat,s323gat);
  nand x74(s376gat,s324gat,s325gat);
  nand x75(s379gat,s326gat,s327gat);
  nand x76(s382gat,s328gat,s329gat);
  nand x77(s385gat,s330gat,s331gat);
  buf x78(s388gat,s290gat);
  buf x79(s389gat,s291gat);
  buf x80(s390gat,s292gat);
  buf x81(s391gat,s297gat);
  or x82(s392gat,s270gat,s343gat);
  not x83(s393gat,s345gat);
  not x84(s399gat,s346gat);
  and x85(s400gat,s348gat,s73gat);
  not x86(s401gat,s349gat);
  not x87(s402gat,s350gat);
  not x88(s403gat,s355gat);
  not x89(s404gat,s357gat);
  not x90(s405gat,s360gat);
  and x91(s406gat,s357gat,s360gat);
  not x92(s407gat,s363gat);
  not x93(s408gat,s366gat);
  and x94(s409gat,s363gat,s366gat);
  nand x95(s410gat,s347gat,s352gat);
  not x96(s411gat,s376gat);
  not x97(s412gat,s379gat);
  and x98(s413gat,s376gat,s379gat);
  not x99(s414gat,s382gat);
  not x100(s415gat,s385gat);
  and x101(s416gat,s382gat,s385gat);
  and x102(s417gat,s210gat,s369gat);
  buf x103(s418gat,s342gat);
  buf x104(s419gat,s344gat);
  buf x105(s420gat,s351gat);
  buf x106(s421gat,s353gat);
  buf x107(s422gat,s354gat);
  buf x108(s423gat,s356gat);
  not x109(s424gat,s400gat);
  and x110(s425gat,s404gat,s405gat);
  and x111(s426gat,s407gat,s408gat);
  and x112(s427gat,s319gat,s393gat,s55gat);
  and x113(s432gat,s393gat,s17gat,s287gat);
  nand x114(s437gat,s393gat,s287gat,s55gat);
  nand x115(s442gat,s375gat,s59gat,s156gat,s393gat);
  nand x116(s443gat,s393gat,s319gat,s17gat);
  and x117(s444gat,s411gat,s412gat);
  and x118(s445gat,s414gat,s415gat);
  buf x119(s446gat,s392gat);
  buf x120(s447gat,s399gat);
  buf x121(s448gat,s401gat);
  buf x122(s449gat,s402gat);
  buf x123(s450gat,s403gat);
  not x124(s451gat,s424gat);
  nor x125(s460gat,s406gat,s425gat);
  nor x126(s463gat,s409gat,s426gat);
  nand x127(s466gat,s442gat,s410gat);
  and x128(s475gat,s143gat,s427gat);
  and x129(s476gat,s310gat,s432gat);
  and x130(s477gat,s146gat,s427gat);
  and x131(s478gat,s310gat,s432gat);
  and x132(s479gat,s149gat,s427gat);
  and x133(s480gat,s310gat,s432gat);
  and x134(s481gat,s153gat,s427gat);
  and x135(s482gat,s310gat,s432gat);
  nand x136(s483gat,s443gat,s1gat);
  or x137(s488gat,s369gat,s437gat);
  or x138(s489gat,s369gat,s437gat);
  or x139(s490gat,s369gat,s437gat);
  or x140(s491gat,s369gat,s437gat);
  nor x141(s492gat,s413gat,s444gat);
  nor x142(s495gat,s416gat,s445gat);
  nand x143(s498gat,s130gat,s460gat);
  or x144(s499gat,s130gat,s460gat);
  nand x145(s500gat,s463gat,s135gat);
  or x146(s501gat,s463gat,s135gat);
  and x147(s502gat,s91gat,s466gat);
  nor x148(s503gat,s475gat,s476gat);
  and x149(s504gat,s96gat,s466gat);
  nor x150(s505gat,s477gat,s478gat);
  and x151(s506gat,s101gat,s466gat);
  nor x152(s507gat,s479gat,s480gat);
  and x153(s508gat,s106gat,s466gat);
  nor x154(s509gat,s481gat,s482gat);
  and x155(s510gat,s143gat,s483gat);
  and x156(s511gat,s111gat,s466gat);
  and x157(s512gat,s146gat,s483gat);
  and x158(s513gat,s116gat,s466gat);
  and x159(s514gat,s149gat,s483gat);
  and x160(s515gat,s121gat,s466gat);
  and x161(s516gat,s153gat,s483gat);
  and x162(s517gat,s126gat,s466gat);
  nand x163(s518gat,s130gat,s492gat);
  or x164(s519gat,s130gat,s492gat);
  nand x165(s520gat,s495gat,s207gat);
  or x166(s521gat,s495gat,s207gat);
  and x167(s522gat,s451gat,s159gat);
  and x168(s523gat,s451gat,s165gat);
  and x169(s524gat,s451gat,s171gat);
  and x170(s525gat,s451gat,s177gat);
  and x171(s526gat,s451gat,s183gat);
  nand x172(s527gat,s451gat,s189gat);
  nand x173(s528gat,s451gat,s195gat);
  nand x174(s529gat,s451gat,s201gat);
  nand x175(s530gat,s498gat,s499gat);
  nand x176(s533gat,s500gat,s501gat);
  nor x177(s536gat,s309gat,s502gat);
  nor x178(s537gat,s316gat,s504gat);
  nor x179(s538gat,s317gat,s506gat);
  nor x180(s539gat,s318gat,s508gat);
  nor x181(s540gat,s510gat,s511gat);
  nor x182(s541gat,s512gat,s513gat);
  nor x183(s542gat,s514gat,s515gat);
  nor x184(s543gat,s516gat,s517gat);
  nand x185(s544gat,s518gat,s519gat);
  nand x186(s547gat,s520gat,s521gat);
  not x187(s550gat,s530gat);
  not x188(s551gat,s533gat);
  and x189(s552gat,s530gat,s533gat);
  nand x190(s553gat,s536gat,s503gat);
  nand x191(s557gat,s537gat,s505gat);
  nand x192(s561gat,s538gat,s507gat);
  nand x193(s565gat,s539gat,s509gat);
  nand x194(s569gat,s488gat,s540gat);
  nand x195(s573gat,s489gat,s541gat);
  nand x196(s577gat,s490gat,s542gat);
  nand x197(s581gat,s491gat,s543gat);
  not x198(s585gat,s544gat);
  not x199(s586gat,s547gat);
  and x200(s587gat,s544gat,s547gat);
  and x201(s588gat,s550gat,s551gat);
  and x202(s589gat,s585gat,s586gat);
  nand x203(s590gat,s553gat,s159gat);
  or x204(s593gat,s553gat,s159gat);
  and x205(s596gat,s246gat,s553gat);
  nand x206(s597gat,s557gat,s165gat);
  or x207(s600gat,s557gat,s165gat);
  and x208(s605gat,s246gat,s557gat);
  nand x209(s606gat,s561gat,s171gat);
  or x210(s609gat,s561gat,s171gat);
  and x211(s615gat,s246gat,s561gat);
  nand x212(s616gat,s565gat,s177gat);
  or x213(s619gat,s565gat,s177gat);
  and x214(s624gat,s246gat,s565gat);
  nand x215(s625gat,s569gat,s183gat);
  or x216(s628gat,s569gat,s183gat);
  and x217(s631gat,s246gat,s569gat);
  nand x218(s632gat,s573gat,s189gat);
  or x219(s635gat,s573gat,s189gat);
  and x220(s640gat,s246gat,s573gat);
  nand x221(s641gat,s577gat,s195gat);
  or x222(s644gat,s577gat,s195gat);
  and x223(s650gat,s246gat,s577gat);
  nand x224(s651gat,s581gat,s201gat);
  or x225(s654gat,s581gat,s201gat);
  and x226(s659gat,s246gat,s581gat);
  nor x227(s660gat,s552gat,s588gat);
  nor x228(s661gat,s587gat,s589gat);
  not x229(s662gat,s590gat);
  and x230(s665gat,s593gat,s590gat);
  nor x231(s669gat,s596gat,s522gat);
  not x232(s670gat,s597gat);
  and x233(s673gat,s600gat,s597gat);
  nor x234(s677gat,s605gat,s523gat);
  not x235(s678gat,s606gat);
  and x236(s682gat,s609gat,s606gat);
  nor x237(s686gat,s615gat,s524gat);
  not x238(s687gat,s616gat);
  and x239(s692gat,s619gat,s616gat);
  nor x240(s696gat,s624gat,s525gat);
  not x241(s697gat,s625gat);
  and x242(s700gat,s628gat,s625gat);
  nor x243(s704gat,s631gat,s526gat);
  not x244(s705gat,s632gat);
  and x245(s708gat,s635gat,s632gat);
  nor x246(s712gat,s337gat,s640gat);
  not x247(s713gat,s641gat);
  and x248(s717gat,s644gat,s641gat);
  nor x249(s721gat,s339gat,s650gat);
  not x250(s722gat,s651gat);
  and x251(s727gat,s654gat,s651gat);
  nor x252(s731gat,s341gat,s659gat);
  nand x253(s732gat,s654gat,s261gat);
  nand x254(s733gat,s644gat,s654gat,s261gat);
  nand x255(s734gat,s635gat,s644gat,s654gat,s261gat);
  not x256(s735gat,s662gat);
  and x257(s736gat,s228gat,s665gat);
  and x258(s737gat,s237gat,s662gat);
  not x259(s738gat,s670gat);
  and x260(s739gat,s228gat,s673gat);
  and x261(s740gat,s237gat,s670gat);
  not x262(s741gat,s678gat);
  and x263(s742gat,s228gat,s682gat);
  and x264(s743gat,s237gat,s678gat);
  not x265(s744gat,s687gat);
  and x266(s745gat,s228gat,s692gat);
  and x267(s746gat,s237gat,s687gat);
  not x268(s747gat,s697gat);
  and x269(s748gat,s228gat,s700gat);
  and x270(s749gat,s237gat,s697gat);
  not x271(s750gat,s705gat);
  and x272(s751gat,s228gat,s708gat);
  and x273(s752gat,s237gat,s705gat);
  not x274(s753gat,s713gat);
  and x275(s754gat,s228gat,s717gat);
  and x276(s755gat,s237gat,s713gat);
  not x277(s756gat,s722gat);
  nor x278(s757gat,s727gat,s261gat);
  and x279(s758gat,s727gat,s261gat);
  and x280(s759gat,s228gat,s727gat);
  and x281(s760gat,s237gat,s722gat);
  nand x282(s761gat,s644gat,s722gat);
  nand x283(s762gat,s635gat,s713gat);
  nand x284(s763gat,s635gat,s644gat,s722gat);
  nand x285(s764gat,s609gat,s687gat);
  nand x286(s765gat,s600gat,s678gat);
  nand x287(s766gat,s600gat,s609gat,s687gat);
  buf x288(s767gat,s660gat);
  buf x289(s768gat,s661gat);
  nor x290(s769gat,s736gat,s737gat);
  nor x291(s770gat,s739gat,s740gat);
  nor x292(s771gat,s742gat,s743gat);
  nor x293(s772gat,s745gat,s746gat);
  nand x294(s773gat,s750gat,s762gat,s763gat,s734gat);
  nor x295(s777gat,s748gat,s749gat);
  nand x296(s778gat,s753gat,s761gat,s733gat);
  nor x297(s781gat,s751gat,s752gat);
  nand x298(s782gat,s756gat,s732gat);
  nor x299(s785gat,s754gat,s755gat);
  nor x300(s786gat,s757gat,s758gat);
  nor x301(s787gat,s759gat,s760gat);
  nor x302(s788gat,s700gat,s773gat);
  and x303(s789gat,s700gat,s773gat);
  nor x304(s790gat,s708gat,s778gat);
  and x305(s791gat,s708gat,s778gat);
  nor x306(s792gat,s717gat,s782gat);
  and x307(s793gat,s717gat,s782gat);
  and x308(s794gat,s219gat,s786gat);
  nand x309(s795gat,s628gat,s773gat);
  nand x310(s796gat,s795gat,s747gat);
  nor x311(s802gat,s788gat,s789gat);
  nor x312(s803gat,s790gat,s791gat);
  nor x313(s804gat,s792gat,s793gat);
  nor x314(s805gat,s340gat,s794gat);
  nor x315(s806gat,s692gat,s796gat);
  and x316(s807gat,s692gat,s796gat);
  and x317(s808gat,s219gat,s802gat);
  and x318(s809gat,s219gat,s803gat);
  and x319(s810gat,s219gat,s804gat);
  nand x320(s811gat,s805gat,s787gat,s731gat,s529gat);
  nand x321(s812gat,s619gat,s796gat);
  nand x322(s813gat,s609gat,s619gat,s796gat);
  nand x323(s814gat,s600gat,s609gat,s619gat,s796gat);
  nand x324(s815gat,s738gat,s765gat,s766gat,s814gat);
  nand x325(s819gat,s741gat,s764gat,s813gat);
  nand x326(s822gat,s744gat,s812gat);
  nor x327(s825gat,s806gat,s807gat);
  nor x328(s826gat,s335gat,s808gat);
  nor x329(s827gat,s336gat,s809gat);
  nor x330(s828gat,s338gat,s810gat);
  not x331(s829gat,s811gat);
  nor x332(s830gat,s665gat,s815gat);
  and x333(s831gat,s665gat,s815gat);
  nor x334(s832gat,s673gat,s819gat);
  and x335(s833gat,s673gat,s819gat);
  nor x336(s834gat,s682gat,s822gat);
  and x337(s835gat,s682gat,s822gat);
  and x338(s836gat,s219gat,s825gat);
  nand x339(s837gat,s826gat,s777gat,s704gat);
  nand x340(s838gat,s827gat,s781gat,s712gat,s527gat);
  nand x341(s839gat,s828gat,s785gat,s721gat,s528gat);
  not x342(s840gat,s829gat);
  nand x343(s841gat,s815gat,s593gat);
  nor x344(s842gat,s830gat,s831gat);
  nor x345(s843gat,s832gat,s833gat);
  nor x346(s844gat,s834gat,s835gat);
  nor x347(s845gat,s334gat,s836gat);
  not x348(s846gat,s837gat);
  not x349(s847gat,s838gat);
  not x350(s848gat,s839gat);
  and x351(s849gat,s735gat,s841gat);
  buf x352(s850gat,s840gat);
  and x353(s851gat,s219gat,s842gat);
  and x354(s852gat,s219gat,s843gat);
  and x355(s853gat,s219gat,s844gat);
  nand x356(s854gat,s845gat,s772gat,s696gat);
  not x357(s855gat,s846gat);
  not x358(s856gat,s847gat);
  not x359(s857gat,s848gat);
  not x360(s858gat,s849gat);
  nor x361(s859gat,s417gat,s851gat);
  nor x362(s860gat,s332gat,s852gat);
  nor x363(s861gat,s333gat,s853gat);
  not x364(s862gat,s854gat);
  buf x365(s863gat,s855gat);
  buf x366(s864gat,s856gat);
  buf x367(s865gat,s857gat);
  buf x368(s866gat,s858gat);
  nand x369(s867gat,s859gat,s769gat,s669gat);
  nand x370(s868gat,s860gat,s770gat,s677gat);
  nand x371(s869gat,s861gat,s771gat,s686gat);
  not x372(s870gat,s862gat);
  not x373(s871gat,s867gat);
  not x374(s872gat,s868gat);
  not x375(s873gat,s869gat);
  buf x376(s874gat,s870gat);
  not x377(s875gat,s871gat);
  not x378(s876gat,s872gat);
  not x379(s877gat,s873gat);
  buf x380(s878gat,s875gat);
  buf x381(s879gat,s876gat);
  buf x382(s880gat,s877gat);

endmodule
