module c7552(s339,s2,s3,s450,s448,s444,s442,s440,s438,s496,s494,s492,s490,s488,s486,s484,s482,s480,s560,s542,s558,s556,s554,s552,s550,s548,s546,s544,s540,s538,s536,s534,s532,s530,s528,s526,s524,s279,s436,s478,s522,s402,s404,s406,s408,s410,s432,s446,s284,s286,s289,s292,s341,s281,s453,s278,s373,s246,s258,s264,s270,s388,s391,s394,s397,s376,s379,s382,s385,s412,s414,s416,s249,s295,s324,s252,s276,s310,s313,s316,s319,s327,s330,s333,s336,s418,s273,s298,s301,s304,s307,s344,s422,s469,s419,s471,s359,s362,s365,s368,s347,s350,s353,s356,s321,s338,s370,s399,s1,s5,s9,s12,s15,s18,s23,s26,s29,s32,s35,s38,s41,s44,s47,s50,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62,s63,s64,s65,s66,s69,s70,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s94,s97,s100,s103,s106,s109,s110,s111,s112,s113,s114,s115,s118,s121,s124,s127,s130,s133,s134,s135,s138,s141,s144,s147,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,s1197,s1455,s1459,s1462,s1469,s1480,s1486,s1492,s1496,s2204,s2208,s2211,s2218,s2224,s2230,s2236,s2239,s2247,s2253,s2256,s3698,s3701,s3705,s3711,s3717,s3723,s3729,s3737,s3743,s3749,s4393,s4394,s4400,s4405,s4410,s4415,s4420,s4427,s4432,s4437,s4526,s4528);

  inout s339;
  output s2;
  output s3;
  output s450;
  output s448;
  output s444;
  output s442;
  output s440;
  output s438;
  output s496;
  output s494;
  output s492;
  output s490;
  output s488;
  output s486;
  output s484;
  output s482;
  output s480;
  output s560;
  output s542;
  output s558;
  output s556;
  output s554;
  output s552;
  output s550;
  output s548;
  output s546;
  output s544;
  output s540;
  output s538;
  output s536;
  output s534;
  output s532;
  output s530;
  output s528;
  output s526;
  output s524;
  output s279;
  output s436;
  output s478;
  output s522;
  output s402;
  output s404;
  output s406;
  output s408;
  output s410;
  output s432;
  output s446;
  output s284;
  output s286;
  output s289;
  output s292;
  output s341;
  output s281;
  output s453;
  output s278;
  output s373;
  output s246;
  output s258;
  output s264;
  output s270;
  output s388;
  output s391;
  output s394;
  output s397;
  output s376;
  output s379;
  output s382;
  output s385;
  output s412;
  output s414;
  output s416;
  output s249;
  output s295;
  output s324;
  output s252;
  output s276;
  output s310;
  output s313;
  output s316;
  output s319;
  output s327;
  output s330;
  output s333;
  output s336;
  output s418;
  output s273;
  output s298;
  output s301;
  output s304;
  output s307;
  output s344;
  output s422;
  output s469;
  output s419;
  output s471;
  output s359;
  output s362;
  output s365;
  output s368;
  output s347;
  output s350;
  output s353;
  output s356;
  output s321;
  output s338;
  output s370;
  output s399;
  input s1;
  input s5;
  input s9;
  input s12;
  input s15;
  input s18;
  input s23;
  input s26;
  input s29;
  input s32;
  input s35;
  input s38;
  input s41;
  input s44;
  input s47;
  input s50;
  input s53;
  input s54;
  input s55;
  input s56;
  input s57;
  input s58;
  input s59;
  input s60;
  input s61;
  input s62;
  input s63;
  input s64;
  input s65;
  input s66;
  input s69;
  input s70;
  input s73;
  input s74;
  input s75;
  input s76;
  input s77;
  input s78;
  input s79;
  input s80;
  input s81;
  input s82;
  input s83;
  input s84;
  input s85;
  input s86;
  input s87;
  input s88;
  input s89;
  input s94;
  input s97;
  input s100;
  input s103;
  input s106;
  input s109;
  input s110;
  input s111;
  input s112;
  input s113;
  input s114;
  input s115;
  input s118;
  input s121;
  input s124;
  input s127;
  input s130;
  input s133;
  input s134;
  input s135;
  input s138;
  input s141;
  input s144;
  input s147;
  input s150;
  input s151;
  input s152;
  input s153;
  input s154;
  input s155;
  input s156;
  input s157;
  input s158;
  input s159;
  input s160;
  input s161;
  input s162;
  input s163;
  input s164;
  input s165;
  input s166;
  input s167;
  input s168;
  input s169;
  input s170;
  input s171;
  input s172;
  input s173;
  input s174;
  input s175;
  input s176;
  input s177;
  input s178;
  input s179;
  input s180;
  input s181;
  input s182;
  input s183;
  input s184;
  input s185;
  input s186;
  input s187;
  input s188;
  input s189;
  input s190;
  input s191;
  input s192;
  input s193;
  input s194;
  input s195;
  input s196;
  input s197;
  input s198;
  input s199;
  input s200;
  input s201;
  input s202;
  input s203;
  input s204;
  input s205;
  input s206;
  input s207;
  input s208;
  input s209;
  input s210;
  input s211;
  input s212;
  input s213;
  input s214;
  input s215;
  input s216;
  input s217;
  input s218;
  input s219;
  input s220;
  input s221;
  input s222;
  input s223;
  input s224;
  input s225;
  input s226;
  input s227;
  input s228;
  input s229;
  input s230;
  input s231;
  input s232;
  input s233;
  input s234;
  input s235;
  input s236;
  input s237;
  input s238;
  input s239;
  input s240;
  input s1197;
  input s1455;
  input s1459;
  input s1462;
  input s1469;
  input s1480;
  input s1486;
  input s1492;
  input s1496;
  input s2204;
  input s2208;
  input s2211;
  input s2218;
  input s2224;
  input s2230;
  input s2236;
  input s2239;
  input s2247;
  input s2253;
  input s2256;
  input s3698;
  input s3701;
  input s3705;
  input s3711;
  input s3717;
  input s3723;
  input s3729;
  input s3737;
  input s3743;
  input s3749;
  input s4393;
  input s4394;
  input s4400;
  input s4405;
  input s4410;
  input s4415;
  input s4420;
  input s4427;
  input s4432;
  input s4437;
  input s4526;
  input s4528;

  buf x0(s2,s1);
  buf x1(s3,s1);
  not x2(s400,s57);
  and x3(s1184,s134,s133);
  buf x4(s450,s1459);
  buf x5(s448,s1469);
  buf x6(s444,s1480);
  buf x7(s442,s1486);
  buf x8(s440,s1492);
  buf x9(s438,s1496);
  and x10(s1501,s162,s172,s188,s199);
  buf x11(s496,s2208);
  buf x12(s494,s2218);
  buf x13(s492,s2224);
  buf x14(s490,s2230);
  buf x15(s488,s2236);
  buf x16(s486,s2239);
  buf x17(s484,s2247);
  buf x18(s482,s2253);
  buf x19(s480,s2256);
  and x20(s2857,s150,s184,s228,s240);
  buf x21(s560,s3698);
  buf x22(s542,s3701);
  buf x23(s558,s3705);
  buf x24(s556,s3711);
  buf x25(s554,s3717);
  buf x26(s552,s3723);
  buf x27(s550,s3729);
  buf x28(s548,s3737);
  buf x29(s546,s3743);
  buf x30(s544,s3749);
  buf x31(s540,s4393);
  buf x32(s538,s4400);
  buf x33(s536,s4405);
  buf x34(s534,s4410);
  buf x35(s532,s4415);
  buf x36(s530,s4420);
  buf x37(s528,s4427);
  buf x38(s526,s4432);
  buf x39(s524,s4437);
  and x40(s4442,s183,s182,s185,s186);
  and x41(s4514,s210,s152,s218,s230);
  not x42(s279,s15);
  not x43(s401,s5);
  buf x44(s573,s1);
  not x45(s574,s5);
  not x46(s575,s5);
  not x47(s1178,s2236);
  not x48(s1186,s2253);
  not x49(s1192,s2256);
  buf x50(s1198,s38);
  buf x51(s1205,s15);
  nand x52(s1206,s12,s9);
  nand x53(s1207,s12,s9);
  buf x54(s1210,s38);
  not x55(s1458,s1455);
  not x56(s1461,s1459);
  buf x57(s436,s1462);
  not x58(s1464,s1462);
  not x59(s1471,s1469);
  buf x60(s1475,s106);
  not x61(s1482,s1480);
  not x62(s1488,s1486);
  not x63(s1495,s1492);
  not x64(s1499,s1496);
  not x65(s1500,s106);
  buf x66(s1503,s18);
  buf x67(s1512,s18);
  and x68(s1518,s4528,s1492);
  buf x69(s1524,s18);
  not x70(s1535,s18);
  nand x71(s1541,s4528,s1496);
  not x72(s2207,s2204);
  not x73(s2210,s2208);
  buf x74(s478,s2211);
  not x75(s2213,s2211);
  not x76(s2220,s2218);
  not x77(s2226,s2224);
  not x78(s2232,s2230);
  not x79(s2238,s2236);
  not x80(s2241,s2239);
  not x81(s2249,s2247);
  not x82(s2255,s2253);
  not x83(s2258,s2256);
  buf x84(s2828,s4526);
  not x85(s3700,s3698);
  not x86(s3703,s3701);
  not x87(s3707,s3705);
  not x88(s3713,s3711);
  not x89(s3719,s3717);
  not x90(s3725,s3723);
  not x91(s3731,s3729);
  not x92(s3739,s3737);
  not x93(s3745,s3743);
  not x94(s3751,s3749);
  not x95(s4121,s4393);
  buf x96(s522,s4394);
  not x97(s4396,s4394);
  not x98(s4402,s4400);
  not x99(s4407,s4405);
  not x100(s4412,s4410);
  not x101(s4417,s4415);
  not x102(s4422,s4420);
  not x103(s4429,s4427);
  not x104(s4434,s4432);
  not x105(s4439,s4437);
  buf x106(s4833,s4526);
  nand x107(s402,s400,s401);
  not x108(s404,s2857);
  not x109(s406,s4514);
  not x110(s408,s4442);
  not x111(s410,s1501);
  and x112(s2876,s2857,s4514);
  and x113(s2878,s4442,s1501);
  buf x114(s432,s573);
  buf x115(s446,s1475);
  not x116(s1519,s1518);
  and x117(s2871,s4528,s1458);
  nand x118(s2883,s4528,s2207);
  and x119(s280,s1184,s575);
  nand x120(s284,s1197,s574);
  not x121(s286,s1205);
  nand x122(s289,s1197,s574);
  nand x123(s292,s1184,s575);
  not x124(s341,s1205);
  not x125(s4839,s4833);
  buf x126(s572,s573);
  buf x127(s581,s1206);
  buf x128(s587,s1512);
  buf x129(s601,s1206);
  buf x130(s606,s1512);
  buf x131(s650,s1206);
  buf x132(s657,s1512);
  buf x133(s671,s1207);
  buf x134(s678,s1503);
  and x135(s777,s1541,s1198);
  and x136(s1115,s1541,s1198);
  buf x137(s1336,s1512);
  buf x138(s1350,s1503);
  not x139(s1477,s1475);
  not x140(s1507,s1503);
  not x141(s1514,s1512);
  not x142(s1530,s1524);
  buf x143(s2259,s1535);
  not x144(s2833,s2828);
  not x145(s2872,s2871);
  buf x146(s2886,s1207);
  buf x147(s2892,s1503);
  buf x148(s2905,s1207);
  buf x149(s2909,s1503);
  buf x150(s3622,s1524);
  buf x151(s3635,s1524);
  buf x152(s3755,s1535);
  buf x153(s4640,s1524);
  buf x154(s4653,s1524);
  buf x155(s4873,s1541);
  buf x156(s4876,s1198);
  buf x157(s4881,s1488);
  buf x158(s4889,s1482);
  buf x159(s4905,s1471);
  buf x160(s4916,s1198);
  buf x161(s4921,s1464);
  buf x162(s5175,s1541);
  buf x163(s5178,s1198);
  buf x164(s5186,s1198);
  buf x165(s5191,s1488);
  buf x166(s5199,s1482);
  buf x167(s5215,s1471);
  buf x168(s5223,s1464);
  buf x169(s5393,s1192);
  buf x170(s5401,s1186);
  buf x171(s5409,s2249);
  buf x172(s5417,s1178);
  buf x173(s5425,s2232);
  buf x174(s5433,s2226);
  buf x175(s5441,s2220);
  buf x176(s5449,s2241);
  buf x177(s5457,s2213);
  buf x178(s5745,s1192);
  buf x179(s5753,s1186);
  buf x180(s5761,s2249);
  buf x181(s5769,s2241);
  buf x182(s5777,s1178);
  buf x183(s5785,s2232);
  buf x184(s5793,s2226);
  buf x185(s5801,s2220);
  buf x186(s5809,s2213);
  buf x187(s5865,s3751);
  buf x188(s5873,s3745);
  buf x189(s5881,s3739);
  buf x190(s5889,s3731);
  buf x191(s5897,s3725);
  buf x192(s5905,s3719);
  buf x193(s5913,s3713);
  buf x194(s5921,s3707);
  buf x195(s5985,s3751);
  buf x196(s5993,s3745);
  buf x197(s6001,s3739);
  buf x198(s6009,s3725);
  buf x199(s6017,s3719);
  buf x200(s6025,s3713);
  buf x201(s6033,s3707);
  buf x202(s6041,s3731);
  buf x203(s6514,s1210);
  buf x204(s6554,s1210);
  buf x205(s6567,s4439);
  buf x206(s6575,s4434);
  buf x207(s6583,s4429);
  buf x208(s6591,s4422);
  buf x209(s6599,s4417);
  buf x210(s6607,s4412);
  buf x211(s6615,s4407);
  buf x212(s6623,s4402);
  buf x213(s6631,s4396);
  buf x214(s6853,s4439);
  buf x215(s6861,s4434);
  buf x216(s6869,s4429);
  buf x217(s6877,s4417);
  buf x218(s6885,s4412);
  buf x219(s6893,s4407);
  buf x220(s6901,s4402);
  buf x221(s6909,s4422);
  buf x222(s6917,s4396);
  not x223(s281,s280);
  buf x224(s453,s572);
  and x225(s784,s1519,s1198);
  and x226(s1014,s1198,s1519);
  and x227(s3221,s2883,s1210);
  buf x228(s4913,s1519);
  nor x229(s4929,s1519,s1198);
  buf x230(s5183,s1519);
  nor x231(s5231,s1198,s1519);
  buf x232(s6511,s2883);
  and x233(s278,s163,s572);
  and x234(s615,s170,s587);
  not x235(s594,s587);
  not x236(s611,s606);
  and x237(s617,s169,s587);
  and x238(s619,s168,s587);
  and x239(s621,s167,s587);
  and x240(s623,s166,s606);
  and x241(s625,s165,s606);
  and x242(s627,s164,s606);
  not x243(s664,s657);
  not x244(s685,s678);
  and x245(s691,s177,s657);
  and x246(s693,s176,s657);
  and x247(s695,s175,s657);
  and x248(s697,s174,s657);
  and x249(s699,s173,s657);
  and x250(s701,s157,s678);
  and x251(s703,s156,s678);
  and x252(s705,s155,s678);
  and x253(s707,s154,s678);
  and x254(s709,s153,s678);
  not x255(s4879,s4873);
  not x256(s4880,s4876);
  not x257(s4887,s4881);
  not x258(s4895,s4889);
  not x259(s4911,s4905);
  not x260(s4920,s4916);
  not x261(s4927,s4921);
  not x262(s5181,s5175);
  not x263(s5182,s5178);
  not x264(s5190,s5186);
  not x265(s5197,s5191);
  not x266(s5205,s5199);
  not x267(s5221,s5215);
  not x268(s5229,s5223);
  not x269(s1343,s1336);
  not x270(s1357,s1350);
  and x271(s1364,s181,s1336);
  and x272(s1366,s171,s1336);
  and x273(s1368,s180,s1336);
  and x274(s1370,s179,s1336);
  and x275(s1372,s178,s1336);
  and x276(s1374,s161,s1350);
  and x277(s1376,s151,s1350);
  and x278(s1378,s160,s1350);
  and x279(s1380,s159,s1350);
  and x280(s1382,s158,s1350);
  not x281(s5399,s5393);
  not x282(s5407,s5401);
  not x283(s5415,s5409);
  not x284(s5423,s5417);
  not x285(s5431,s5425);
  not x286(s5439,s5433);
  not x287(s5447,s5441);
  not x288(s5455,s5449);
  not x289(s5463,s5457);
  not x290(s5751,s5745);
  not x291(s5759,s5753);
  not x292(s5767,s5761);
  not x293(s5775,s5769);
  not x294(s5783,s5777);
  not x295(s5791,s5785);
  not x296(s5799,s5793);
  not x297(s5807,s5801);
  not x298(s5815,s5809);
  buf x299(s2019,s1514);
  buf x300(s2032,s1507);
  buf x301(s2117,s1514);
  buf x302(s2130,s1507);
  not x303(s2266,s2259);
  buf x304(s2272,s1507);
  and x305(s2286,s44,s2259);
  and x306(s2288,s41,s2259);
  and x307(s2290,s29,s2259);
  and x308(s2292,s26,s2259);
  and x309(s2294,s23,s2259);
  not x310(s5871,s5865);
  not x311(s5879,s5873);
  not x312(s5887,s5881);
  not x313(s5895,s5889);
  not x314(s5903,s5897);
  not x315(s5911,s5905);
  not x316(s5919,s5913);
  not x317(s5927,s5921);
  not x318(s5991,s5985);
  not x319(s5999,s5993);
  not x320(s6007,s6001);
  not x321(s6015,s6009);
  not x322(s6023,s6017);
  not x323(s6031,s6025);
  not x324(s6039,s6033);
  not x325(s6047,s6041);
  not x326(s2899,s2892);
  not x327(s2914,s2909);
  and x328(s2919,s209,s2892);
  and x329(s2921,s216,s2892);
  and x330(s2923,s215,s2892);
  and x331(s2925,s214,s2892);
  and x332(s2927,s213,s2909);
  and x333(s2929,s212,s2909);
  and x334(s2931,s211,s2909);
  not x335(s6518,s6514);
  and x336(s3173,s2872,s1210);
  not x337(s6558,s6554);
  not x338(s6573,s6567);
  not x339(s6581,s6575);
  not x340(s6589,s6583);
  not x341(s6597,s6591);
  not x342(s6605,s6599);
  not x343(s6613,s6607);
  not x344(s6621,s6615);
  not x345(s6629,s6623);
  not x346(s6637,s6631);
  not x347(s3629,s3622);
  not x348(s3642,s3635);
  and x349(s3649,s1461,s3622);
  and x350(s3651,s1464,s3622);
  and x351(s3653,s1471,s3622);
  and x352(s3655,s1500,s3622);
  and x353(s3657,s1482,s3622);
  and x354(s3659,s1488,s3635);
  and x355(s3661,s1495,s3635);
  and x356(s3663,s1499,s3635);
  not x357(s3762,s3755);
  buf x358(s3768,s1507);
  and x359(s3782,s47,s3755);
  and x360(s3784,s35,s3755);
  and x361(s3786,s32,s3755);
  and x362(s3788,s50,s3755);
  and x363(s3790,s66,s3755);
  not x364(s6859,s6853);
  not x365(s6867,s6861);
  not x366(s6875,s6869);
  not x367(s6883,s6877);
  not x368(s6891,s6885);
  not x369(s6899,s6893);
  not x370(s6907,s6901);
  not x371(s6915,s6909);
  not x372(s6923,s6917);
  buf x373(s4094,s1530);
  buf x374(s4107,s1530);
  buf x375(s4444,s1530);
  buf x376(s4457,s1530);
  not x377(s4647,s4640);
  not x378(s4660,s4653);
  and x379(s4667,s2210,s4640);
  and x380(s4669,s2213,s4640);
  and x381(s4671,s2220,s4640);
  and x382(s4673,s2226,s4640);
  and x383(s4675,s2232,s4640);
  and x384(s4677,s2238,s4653);
  and x385(s4679,s2241,s4653);
  and x386(s4681,s2249,s4653);
  and x387(s4683,s2255,s4653);
  and x388(s4685,s2258,s4653);
  buf x389(s4897,s1477);
  buf x390(s5207,s1477);
  buf x391(s6551,s2872);
  nand x392(s763,s4876,s4879);
  nand x393(s764,s4873,s4880);
  not x394(s4919,s4913);
  nand x395(s886,s4913,s4920);
  nand x396(s1005,s5178,s5181);
  nand x397(s1006,s5175,s5182);
  not x398(s5189,s5183);
  nand x399(s1018,s5183,s5190);
  not x400(s5237,s5231);
  not x401(s6517,s6511);
  nand x402(s3169,s6511,s6518);
  not x403(s4935,s4929);
  buf x404(s4970,s784);
  buf x405(s5239,s1014);
  or x406(s577,s594,s615);
  or x407(s616,s594,s587);
  or x408(s618,s594,s617);
  or x409(s620,s594,s619);
  or x410(s622,s594,s621);
  or x411(s624,s611,s623);
  or x412(s626,s611,s625);
  or x413(s628,s611,s627);
  or x414(s692,s664,s691);
  or x415(s694,s664,s693);
  or x416(s696,s664,s695);
  or x417(s698,s664,s697);
  or x418(s700,s664,s699);
  or x419(s702,s685,s701);
  or x420(s704,s685,s703);
  or x421(s706,s685,s705);
  or x422(s708,s685,s707);
  or x423(s710,s685,s709);
  nand x424(s765,s763,s764);
  not x425(s4903,s4897);
  nand x426(s885,s4916,s4919);
  nand x427(s1007,s1005,s1006);
  nand x428(s1017,s5186,s5189);
  not x429(s5213,s5207);
  and x430(s1363,s141,s1343);
  and x431(s1365,s147,s1343);
  and x432(s1367,s138,s1343);
  and x433(s1369,s144,s1343);
  and x434(s1371,s135,s1343);
  and x435(s1373,s141,s1357);
  and x436(s1375,s147,s1357);
  and x437(s1377,s138,s1357);
  and x438(s1379,s144,s1357);
  and x439(s1381,s135,s1357);
  not x440(s2026,s2019);
  not x441(s2039,s2032);
  and x442(s2046,s103,s2019);
  and x443(s2048,s130,s2019);
  and x444(s2050,s127,s2019);
  and x445(s2052,s124,s2019);
  and x446(s2054,s100,s2019);
  and x447(s2056,s103,s2032);
  and x448(s2058,s130,s2032);
  and x449(s2060,s127,s2032);
  and x450(s2062,s124,s2032);
  and x451(s2064,s100,s2032);
  not x452(s2124,s2117);
  not x453(s2137,s2130);
  and x454(s2144,s115,s2117);
  and x455(s2146,s118,s2117);
  and x456(s2148,s97,s2117);
  and x457(s2150,s94,s2117);
  and x458(s2152,s121,s2117);
  and x459(s2154,s115,s2130);
  and x460(s2156,s118,s2130);
  and x461(s2158,s97,s2130);
  and x462(s2160,s94,s2130);
  and x463(s2162,s121,s2130);
  not x464(s2279,s2272);
  and x465(s2285,s208,s2266);
  and x466(s2287,s198,s2266);
  and x467(s2289,s207,s2266);
  and x468(s2291,s206,s2266);
  and x469(s2293,s205,s2266);
  and x470(s2296,s44,s2272);
  and x471(s2298,s41,s2272);
  and x472(s2300,s29,s2272);
  and x473(s2302,s26,s2272);
  and x474(s2304,s23,s2272);
  or x475(s2918,s2899,s2892);
  or x476(s2920,s2899,s2919);
  or x477(s2922,s2899,s2921);
  or x478(s2924,s2899,s2923);
  or x479(s2926,s2899,s2925);
  or x480(s2928,s2914,s2927);
  or x481(s2930,s2914,s2929);
  or x482(s2932,s2914,s2931);
  nand x483(s3168,s6514,s6517);
  not x484(s6557,s6551);
  nand x485(s3211,s6551,s6558);
  and x486(s3648,s114,s3629);
  and x487(s3650,s113,s3629);
  and x488(s3652,s111,s3629);
  and x489(s3654,s87,s3629);
  and x490(s3656,s112,s3629);
  and x491(s3658,s88,s3642);
  and x492(s3660,s1455,s3642);
  and x493(s3662,s2204,s3642);
  and x494(s3665,s3703,s3642);
  and x495(s3666,s70,s3642);
  not x496(s3775,s3768);
  and x497(s3781,s193,s3762);
  and x498(s3783,s192,s3762);
  and x499(s3785,s191,s3762);
  and x500(s3787,s190,s3762);
  and x501(s3789,s189,s3762);
  and x502(s3792,s47,s3768);
  and x503(s3794,s35,s3768);
  and x504(s3796,s32,s3768);
  and x505(s3798,s50,s3768);
  and x506(s3800,s66,s3768);
  not x507(s4101,s4094);
  not x508(s4114,s4107);
  and x509(s4123,s58,s4094);
  and x510(s4126,s77,s4094);
  and x511(s4129,s78,s4094);
  and x512(s4132,s59,s4094);
  and x513(s4135,s81,s4094);
  and x514(s4138,s80,s4107);
  and x515(s4141,s79,s4107);
  and x516(s4144,s60,s4107);
  and x517(s4147,s61,s4107);
  and x518(s4150,s62,s4107);
  not x519(s4451,s4444);
  not x520(s4464,s4457);
  and x521(s4471,s69,s4444);
  and x522(s4473,s70,s4444);
  and x523(s4475,s74,s4444);
  and x524(s4477,s76,s4444);
  and x525(s4479,s75,s4444);
  and x526(s4481,s73,s4457);
  and x527(s4483,s53,s4457);
  and x528(s4485,s54,s4457);
  and x529(s4487,s55,s4457);
  and x530(s4489,s56,s4457);
  and x531(s4666,s82,s4647);
  and x532(s4668,s65,s4647);
  and x533(s4670,s83,s4647);
  and x534(s4672,s84,s4647);
  and x535(s4674,s85,s4647);
  and x536(s4676,s64,s4660);
  and x537(s4678,s63,s4660);
  and x538(s4680,s86,s4660);
  and x539(s4682,s109,s4660);
  and x540(s4684,s110,s4660);
  and x541(s579,s577,s581);
  and x542(s629,s616,s581);
  and x543(s633,s618,s581);
  and x544(s637,s620,s581);
  and x545(s641,s622,s581);
  and x546(s645,s624,s601);
  and x547(s711,s692,s650);
  and x548(s715,s694,s650);
  and x549(s719,s696,s650);
  and x550(s723,s698,s650);
  and x551(s727,s700,s650);
  and x552(s731,s702,s671);
  and x553(s737,s704,s671);
  and x554(s745,s706,s671);
  and x555(s751,s708,s671);
  and x556(s757,s710,s671);
  nand x557(s887,s885,s886);
  nand x558(s1019,s1017,s1018);
  not x559(s5245,s5239);
  or x560(s1383,s1365,s1366);
  or x561(s1387,s1367,s1368);
  or x562(s1391,s1369,s1370);
  or x563(s1395,s1371,s1372);
  or x564(s1399,s1375,s1376);
  or x565(s1406,s1377,s1378);
  or x566(s1412,s1379,s1380);
  or x567(s1418,s1381,s1382);
  or x568(s2305,s2287,s2288);
  or x569(s2308,s2289,s2290);
  or x570(s2312,s2291,s2292);
  or x571(s2316,s2293,s2294);
  and x572(s2933,s2920,s2886);
  and x573(s2938,s2922,s2886);
  and x574(s2942,s2924,s2886);
  and x575(s2946,s2926,s2886);
  and x576(s2950,s2928,s2905);
  nand x577(s3170,s3168,s3169);
  nand x578(s3210,s6554,s6557);
  or x579(s3667,s3650,s3651);
  or x580(s3670,s3652,s3653);
  or x581(s3673,s3654,s3655);
  or x582(s3676,s3656,s3657);
  or x583(s3679,s3658,s3659);
  or x584(s3682,s3665,s3635);
  or x585(s3686,s3666,s3635);
  or x586(s3801,s3781,s3782);
  or x587(s3804,s3783,s3784);
  or x588(s3807,s3785,s3786);
  or x589(s3810,s3787,s3788);
  or x590(s3813,s3789,s3790);
  and x591(s4525,s2918,s2886);
  or x592(s4686,s4668,s4669);
  or x593(s4689,s4670,s4671);
  or x594(s4692,s4672,s4673);
  or x595(s4695,s4674,s4675);
  or x596(s4698,s4676,s4677);
  or x597(s4701,s4678,s4679);
  or x598(s4704,s4680,s4681);
  or x599(s4707,s4682,s4683);
  or x600(s4710,s4684,s4685);
  not x601(s4976,s4970);
  and x602(s5271,s2932,s2905);
  and x603(s5274,s2930,s2905);
  and x604(s5305,s628,s601);
  and x605(s5308,s626,s601);
  or x606(s5318,s1373,s1374);
  or x607(s6690,s3648,s3649);
  or x608(s6711,s3662,s3663);
  or x609(s6714,s3660,s3661);
  or x610(s7252,s2285,s2286);
  or x611(s7296,s1363,s1364);
  or x612(s7466,s4666,s4667);
  and x613(s907,s765,s784);
  and x614(s913,s765,s784);
  and x615(s915,s765,s784);
  and x616(s916,s765,s784);
  and x617(s1116,s1007,s1014);
  and x618(s2045,s204,s2026);
  and x619(s2047,s203,s2026);
  and x620(s2049,s202,s2026);
  and x621(s2051,s201,s2026);
  and x622(s2053,s200,s2026);
  and x623(s2055,s235,s2039);
  and x624(s2057,s234,s2039);
  and x625(s2059,s233,s2039);
  and x626(s2061,s232,s2039);
  and x627(s2063,s231,s2039);
  and x628(s2143,s197,s2124);
  and x629(s2145,s187,s2124);
  and x630(s2147,s196,s2124);
  and x631(s2149,s195,s2124);
  and x632(s2151,s194,s2124);
  and x633(s2153,s227,s2137);
  and x634(s2155,s217,s2137);
  and x635(s2157,s226,s2137);
  and x636(s2159,s225,s2137);
  and x637(s2161,s224,s2137);
  and x638(s2295,s239,s2279);
  and x639(s2297,s229,s2279);
  and x640(s2299,s238,s2279);
  and x641(s2301,s237,s2279);
  and x642(s2303,s236,s2279);
  nand x643(s3212,s3210,s3211);
  and x644(s3791,s223,s3775);
  and x645(s3793,s222,s3775);
  and x646(s3795,s221,s3775);
  and x647(s3797,s220,s3775);
  and x648(s3799,s219,s3775);
  and x649(s4122,s4121,s4101);
  and x650(s4125,s4396,s4101);
  and x651(s4128,s4402,s4101);
  and x652(s4131,s4407,s4101);
  and x653(s4134,s4412,s4101);
  and x654(s4137,s4417,s4114);
  and x655(s4140,s4422,s4114);
  and x656(s4143,s4429,s4114);
  and x657(s4146,s4434,s4114);
  and x658(s4149,s4439,s4114);
  and x659(s4470,s3700,s4451);
  and x660(s4472,s3703,s4451);
  and x661(s4474,s3707,s4451);
  and x662(s4476,s3713,s4451);
  and x663(s4478,s3719,s4451);
  and x664(s4480,s3725,s4464);
  and x665(s4482,s3731,s4464);
  and x666(s4484,s3739,s4464);
  and x667(s4486,s3745,s4464);
  and x668(s4488,s3751,s4464);
  buf x669(s4962,s765);
  buf x670(s5003,s765);
  buf x671(s5234,s1007);
  buf x672(s5242,s1007);
  not x673(s5250,s4525);
  not x674(s5284,s579);
  and x675(s802,s1488,s2950);
  and x676(s821,s1482,s2946);
  and x677(s845,s1477,s2942);
  and x678(s868,s1471,s2938);
  and x679(s877,s1464,s2933);
  and x680(s902,s887,s765);
  or x681(s908,s777,s907);
  and x682(s914,s887,s765);
  or x683(s917,s777,s916);
  and x684(s953,s887,s765);
  not x685(s1023,s1019);
  and x686(s1035,s1488,s2950);
  and x687(s1050,s1482,s2946);
  and x688(s1068,s1477,s2942);
  and x689(s1086,s1471,s2938);
  and x690(s1102,s1464,s2933);
  and x691(s1108,s1019,s1007);
  or x692(s1117,s1115,s1116);
  not x693(s5322,s5318);
  and x694(s1553,s1192,s757);
  and x695(s1567,s1186,s751);
  and x696(s1584,s2249,s745);
  and x697(s1590,s2241,s737);
  and x698(s1606,s1178,s731);
  and x699(s1624,s2232,s1418);
  and x700(s1647,s2226,s1412);
  and x701(s1669,s2220,s1406);
  and x702(s1677,s2213,s1399);
  and x703(s1802,s1192,s757);
  and x704(s1816,s1186,s751);
  and x705(s1834,s2249,s745);
  and x706(s1841,s737,s2241);
  and x707(s1866,s1178,s731);
  and x708(s1880,s2232,s1418);
  and x709(s1897,s2226,s1412);
  and x710(s1914,s2220,s1406);
  and x711(s1929,s2213,s1399);
  or x712(s2065,s2045,s2046);
  or x713(s2069,s2047,s2048);
  or x714(s2073,s2049,s2050);
  or x715(s2077,s2051,s2052);
  or x716(s2081,s2053,s2054);
  or x717(s2085,s2055,s2056);
  or x718(s2091,s2057,s2058);
  or x719(s2099,s2059,s2060);
  or x720(s2105,s2061,s2062);
  or x721(s2111,s2063,s2064);
  or x722(s2163,s2145,s2146);
  or x723(s2167,s2147,s2148);
  or x724(s2171,s2149,s2150);
  or x725(s2175,s2151,s2152);
  or x726(s2179,s2155,s2156);
  or x727(s2186,s2157,s2158);
  or x728(s2192,s2159,s2160);
  or x729(s2198,s2161,s2162);
  or x730(s2320,s2297,s2298);
  or x731(s2323,s2299,s2300);
  or x732(s2329,s2301,s2302);
  or x733(s2335,s2303,s2304);
  and x734(s2962,s4710,s727);
  and x735(s2970,s4707,s723);
  and x736(s2977,s4704,s719);
  and x737(s2979,s4701,s715);
  and x738(s2989,s4698,s711);
  and x739(s2998,s4695,s1395);
  and x740(s3006,s4692,s1391);
  and x741(s3013,s4689,s1387);
  and x742(s3015,s4686,s1383);
  and x743(s3183,s3679,s645);
  and x744(s3192,s3676,s641);
  and x745(s3200,s3673,s637);
  and x746(s3207,s3670,s633);
  and x747(s3209,s3667,s629);
  and x748(s3216,s3212,s3170);
  and x749(s3222,s3170,s3173);
  not x750(s6694,s6690);
  and x751(s3695,s1535,s2305);
  or x752(s3816,s3791,s3792);
  or x753(s3821,s3793,s3794);
  or x754(s3828,s3795,s3796);
  or x755(s3833,s3797,s3798);
  or x756(s3838,s3799,s3800);
  or x757(s4151,s4125,s4126);
  or x758(s4154,s4128,s4129);
  or x759(s4157,s4131,s4132);
  or x760(s4160,s4134,s4135);
  or x761(s4163,s4137,s4138);
  or x762(s4166,s4140,s4141);
  or x763(s4169,s4143,s4144);
  or x764(s4172,s4146,s4147);
  or x765(s4175,s4149,s4150);
  not x766(s7256,s7252);
  not x767(s7300,s7296);
  or x768(s4490,s4474,s4475);
  or x769(s4493,s4476,s4477);
  or x770(s4496,s4478,s4479);
  or x771(s4499,s4480,s4481);
  or x772(s4502,s4482,s4483);
  or x773(s4505,s4484,s4485);
  or x774(s4508,s4486,s4487);
  or x775(s4511,s4488,s4489);
  not x776(s7470,s7466);
  buf x777(s4884,s2950);
  buf x778(s4892,s2946);
  buf x779(s4900,s2942);
  buf x780(s4908,s2938);
  buf x781(s4924,s2933);
  buf x782(s4952,s887);
  nor x783(s4983,s777,s915);
  buf x784(s4993,s887);
  nor x785(s5011,s1464,s2933);
  buf x786(s5194,s2950);
  buf x787(s5202,s2946);
  buf x788(s5210,s2942);
  buf x789(s5218,s2938);
  buf x790(s5226,s2933);
  buf x791(s5247,s2933);
  buf x792(s5255,s2942);
  buf x793(s5258,s2938);
  buf x794(s5263,s2950);
  buf x795(s5266,s2946);
  not x796(s5277,s5271);
  not x797(s5278,s5274);
  buf x798(s5281,s629);
  buf x799(s5289,s637);
  buf x800(s5292,s633);
  buf x801(s5297,s645);
  buf x802(s5300,s641);
  not x803(s5311,s5305);
  not x804(s5312,s5308);
  buf x805(s5315,s1399);
  buf x806(s5323,s1412);
  buf x807(s5326,s1406);
  buf x808(s5331,s731);
  buf x809(s5334,s1418);
  buf x810(s5339,s745);
  buf x811(s5342,s737);
  buf x812(s5349,s757);
  buf x813(s5352,s751);
  buf x814(s5396,s757);
  buf x815(s5404,s751);
  buf x816(s5412,s745);
  buf x817(s5420,s731);
  buf x818(s5428,s1418);
  buf x819(s5436,s1412);
  buf x820(s5444,s1406);
  buf x821(s5452,s737);
  buf x822(s5460,s1399);
  nor x823(s5465,s2241,s737);
  nor x824(s5581,s2213,s1399);
  buf x825(s5748,s757);
  buf x826(s5756,s751);
  buf x827(s5764,s745);
  buf x828(s5772,s737);
  buf x829(s5780,s731);
  buf x830(s5788,s1418);
  buf x831(s5796,s1412);
  buf x832(s5804,s1406);
  buf x833(s5812,s1399);
  nor x834(s5849,s737,s2241);
  buf x835(s5929,s3682);
  buf x836(s6049,s3682);
  buf x837(s6367,s4710);
  buf x838(s6370,s727);
  buf x839(s6375,s4707);
  buf x840(s6378,s723);
  buf x841(s6383,s4704);
  buf x842(s6386,s719);
  buf x843(s6391,s4698);
  buf x844(s6394,s711);
  buf x845(s6399,s4695);
  buf x846(s6402,s1395);
  buf x847(s6407,s4692);
  buf x848(s6410,s1391);
  buf x849(s6415,s4689);
  buf x850(s6418,s1387);
  buf x851(s6423,s4701);
  buf x852(s6426,s715);
  buf x853(s6431,s4686);
  buf x854(s6434,s1383);
  buf x855(s6442,s3813);
  buf x856(s6450,s3810);
  buf x857(s6458,s3807);
  buf x858(s6466,s3801);
  buf x859(s6498,s3804);
  buf x860(s6519,s3679);
  buf x861(s6522,s645);
  buf x862(s6527,s3676);
  buf x863(s6530,s641);
  buf x864(s6535,s3673);
  buf x865(s6538,s637);
  buf x866(s6543,s3670);
  buf x867(s6546,s633);
  buf x868(s6559,s3667);
  buf x869(s6562,s629);
  buf x870(s6687,s3667);
  buf x871(s6695,s3673);
  buf x872(s6698,s3670);
  buf x873(s6703,s3679);
  buf x874(s6706,s3676);
  not x875(s6717,s6711);
  not x876(s6718,s6714);
  or x877(s6724,s2153,s2154);
  or x878(s6768,s2295,s2296);
  or x879(s7208,s2143,s2144);
  buf x880(s7221,s3801);
  buf x881(s7229,s3807);
  buf x882(s7232,s3804);
  buf x883(s7239,s3813);
  buf x884(s7242,s3810);
  buf x885(s7249,s2305);
  buf x886(s7257,s2312);
  buf x887(s7260,s2308);
  buf x888(s7268,s2316);
  buf x889(s7293,s1383);
  buf x890(s7301,s1391);
  buf x891(s7304,s1387);
  buf x892(s7309,s711);
  buf x893(s7312,s1395);
  buf x894(s7317,s719);
  buf x895(s7320,s715);
  buf x896(s7327,s727);
  buf x897(s7330,s723);
  buf x898(s7396,s2316);
  buf x899(s7404,s2312);
  buf x900(s7412,s2308);
  buf x901(s7425,s3686);
  buf x902(s7463,s4686);
  buf x903(s7471,s4692);
  buf x904(s7474,s4689);
  buf x905(s7479,s4698);
  buf x906(s7482,s4695);
  buf x907(s7487,s4704);
  buf x908(s7490,s4701);
  buf x909(s7497,s4710);
  buf x910(s7500,s4707);
  or x911(s7507,s4472,s4473);
  or x912(s7510,s4470,s4471);
  or x913(s7554,s4122,s4123);
  nand x914(s1152,s5234,s5237);
  not x915(s5238,s5234);
  nand x916(s1156,s5242,s5245);
  not x917(s5246,s5242);
  not x918(s5254,s5250);
  not x919(s5288,s5284);
  or x920(s3223,s3221,s3222);
  or x921(s4942,s777,s913,s914);
  not x922(s4966,s4962);
  not x923(s5007,s5003);
  nand x924(s5279,s5274,s5277);
  nand x925(s5280,s5271,s5278);
  nand x926(s5313,s5308,s5311);
  nand x927(s5314,s5305,s5312);
  nand x928(s6719,s6714,s6717);
  nand x929(s6720,s6711,s6718);
  nand x930(s790,s4884,s4887);
  not x931(s4888,s4884);
  nand x932(s803,s4892,s4895);
  not x933(s4896,s4892);
  nand x934(s825,s4900,s4903);
  not x935(s4904,s4900);
  nand x936(s851,s4908,s4911);
  not x937(s4912,s4908);
  nand x938(s893,s4924,s4927);
  not x939(s4928,s4924);
  not x940(s906,s902);
  not x941(s912,s908);
  nand x942(s1024,s5194,s5197);
  not x943(s5198,s5194);
  nand x944(s1036,s5202,s5205);
  not x945(s5206,s5202);
  nand x946(s1053,s5210,s5213);
  not x947(s5214,s5210);
  nand x948(s1072,s5218,s5221);
  not x949(s5222,s5218);
  nand x950(s1091,s5226,s5229);
  not x951(s5230,s5226);
  not x952(s1112,s1108);
  not x953(s1121,s1117);
  nand x954(s1153,s5231,s5238);
  nand x955(s1157,s5239,s5246);
  not x956(s5253,s5247);
  nand x957(s1216,s5247,s5254);
  not x958(s5261,s5255);
  not x959(s5262,s5258);
  not x960(s5269,s5263);
  not x961(s5270,s5266);
  not x962(s5287,s5281);
  nand x963(s1239,s5281,s5288);
  not x964(s5295,s5289);
  not x965(s5296,s5292);
  not x966(s5303,s5297);
  not x967(s5304,s5300);
  not x968(s5321,s5315);
  nand x969(s1262,s5315,s5322);
  not x970(s5329,s5323);
  not x971(s5330,s5326);
  not x972(s5337,s5331);
  not x973(s5338,s5334);
  nand x974(s1544,s5396,s5399);
  not x975(s5400,s5396);
  nand x976(s1554,s5404,s5407);
  not x977(s5408,s5404);
  nand x978(s1571,s5412,s5415);
  not x979(s5416,s5412);
  nand x980(s1596,s5420,s5423);
  not x981(s5424,s5420);
  nand x982(s1607,s5428,s5431);
  not x983(s5432,s5428);
  nand x984(s1628,s5436,s5439);
  not x985(s5440,s5436);
  nand x986(s1653,s5444,s5447);
  not x987(s5448,s5444);
  nand x988(s1685,s5452,s5455);
  not x989(s5456,s5452);
  nand x990(s1693,s5460,s5463);
  not x991(s5464,s5460);
  nand x992(s1793,s5748,s5751);
  not x993(s5752,s5748);
  nand x994(s1803,s5756,s5759);
  not x995(s5760,s5756);
  nand x996(s1820,s5764,s5767);
  not x997(s5768,s5764);
  nand x998(s1848,s5772,s5775);
  not x999(s5776,s5772);
  nand x1000(s1857,s5780,s5783);
  not x1001(s5784,s5780);
  nand x1002(s1867,s5788,s5791);
  not x1003(s5792,s5788);
  nand x1004(s1883,s5796,s5799);
  not x1005(s5800,s5796);
  nand x1006(s1901,s5804,s5807);
  not x1007(s5808,s5804);
  nand x1008(s1919,s5812,s5815);
  not x1009(s5816,s5812);
  not x1010(s5855,s5849);
  and x1011(s2351,s3751,s2111);
  and x1012(s2366,s3745,s2105);
  and x1013(s2384,s3739,s2099);
  and x1014(s2391,s2091,s3731);
  and x1015(s2417,s3725,s2085);
  and x1016(s2431,s3719,s2335);
  and x1017(s2448,s3713,s2329);
  and x1018(s2465,s3707,s2323);
  not x1019(s5935,s5929);
  and x1020(s2597,s3751,s2111);
  and x1021(s2612,s3745,s2105);
  and x1022(s2629,s3739,s2099);
  and x1023(s2635,s3731,s2091);
  and x1024(s2652,s3725,s2085);
  and x1025(s2670,s3719,s2335);
  and x1026(s2693,s3713,s2329);
  and x1027(s2715,s3707,s2323);
  not x1028(s6055,s6049);
  not x1029(s6373,s6367);
  not x1030(s6374,s6370);
  not x1031(s6381,s6375);
  not x1032(s6382,s6378);
  not x1033(s6389,s6383);
  not x1034(s6390,s6386);
  not x1035(s6397,s6391);
  not x1036(s6398,s6394);
  not x1037(s6405,s6399);
  not x1038(s6406,s6402);
  not x1039(s6413,s6407);
  not x1040(s6414,s6410);
  not x1041(s6421,s6415);
  not x1042(s6422,s6418);
  not x1043(s6429,s6423);
  not x1044(s6430,s6426);
  not x1045(s6437,s6431);
  not x1046(s6438,s6434);
  not x1047(s6446,s6442);
  and x1048(s3059,s4175,s3813);
  not x1049(s6454,s6450);
  and x1050(s3068,s4172,s3810);
  not x1051(s6462,s6458);
  and x1052(s3076,s4169,s3807);
  and x1053(s3079,s4166,s3804);
  not x1054(s6470,s6466);
  and x1055(s3090,s4163,s3801);
  and x1056(s3099,s4160,s2175);
  and x1057(s3107,s4157,s2171);
  and x1058(s3114,s4154,s2167);
  and x1059(s3116,s4151,s2163);
  not x1060(s6502,s6498);
  not x1061(s6525,s6519);
  not x1062(s6526,s6522);
  not x1063(s6533,s6527);
  not x1064(s6534,s6530);
  not x1065(s6541,s6535);
  not x1066(s6542,s6538);
  not x1067(s6549,s6543);
  not x1068(s6550,s6546);
  not x1069(s6565,s6559);
  not x1070(s6566,s6562);
  not x1071(s3220,s3216);
  and x1072(s3292,s4439,s3838);
  and x1073(s3308,s4434,s3833);
  and x1074(s3327,s4429,s3828);
  and x1075(s3335,s3821,s4422);
  and x1076(s3362,s4417,s3816);
  and x1077(s3376,s4412,s2198);
  and x1078(s3393,s4407,s2192);
  and x1079(s3410,s4402,s2186);
  and x1080(s3425,s4396,s2179);
  not x1081(s6693,s6687);
  nand x1082(s3503,s6687,s6694);
  not x1083(s6701,s6695);
  not x1084(s6702,s6698);
  not x1085(s6709,s6703);
  not x1086(s6710,s6706);
  not x1087(s6728,s6724);
  not x1088(s6772,s6768);
  and x1089(s3853,s4439,s3838);
  and x1090(s3868,s4434,s3833);
  and x1091(s3885,s4429,s3828);
  and x1092(s3891,s4422,s3821);
  and x1093(s3908,s4417,s3816);
  and x1094(s3926,s4412,s2198);
  and x1095(s3949,s4407,s2192);
  and x1096(s3971,s4402,s2186);
  and x1097(s3979,s4396,s2179);
  not x1098(s7212,s7208);
  not x1099(s7227,s7221);
  not x1100(s7255,s7249);
  nand x1101(s4202,s7249,s7256);
  not x1102(s7263,s7257);
  not x1103(s7264,s7260);
  not x1104(s7272,s7268);
  not x1105(s7299,s7293);
  nand x1106(s4225,s7293,s7300);
  not x1107(s7307,s7301);
  not x1108(s7308,s7304);
  not x1109(s7315,s7309);
  not x1110(s7316,s7312);
  and x1111(s4297,s4511,s2081);
  and x1112(s4305,s4508,s2077);
  and x1113(s4312,s4505,s2073);
  and x1114(s4314,s4502,s2069);
  and x1115(s4324,s4499,s2065);
  not x1116(s7400,s7396);
  and x1117(s4333,s4496,s2316);
  not x1118(s7408,s7404);
  and x1119(s4341,s4493,s2312);
  not x1120(s7416,s7412);
  and x1121(s4348,s4490,s2308);
  and x1122(s4349,s3686,s3695);
  not x1123(s7431,s7425);
  and x1124(s4389,s2320,s1535);
  not x1125(s7469,s7463);
  nand x1126(s4530,s7463,s7470);
  not x1127(s7477,s7471);
  not x1128(s7478,s7474);
  not x1129(s7485,s7479);
  not x1130(s7486,s7482);
  not x1131(s7513,s7507);
  not x1132(s7514,s7510);
  not x1133(s7558,s7554);
  or x1134(s4932,s917,s953);
  not x1135(s4956,s4952);
  not x1136(s4973,s917);
  not x1137(s4987,s4983);
  not x1138(s4997,s4993);
  not x1139(s5017,s5011);
  buf x1140(s5099,s877);
  not x1141(s5345,s5339);
  not x1142(s5346,s5342);
  not x1143(s5355,s5349);
  not x1144(s5356,s5352);
  nand x1145(s5372,s5279,s5280);
  nand x1146(s5380,s5313,s5314);
  not x1147(s5471,s5465);
  buf x1148(s5523,s1590);
  not x1149(s5587,s5581);
  buf x1150(s5669,s1677);
  buf x1151(s5857,s1841);
  buf x1152(s5868,s2111);
  buf x1153(s5876,s2105);
  buf x1154(s5884,s2099);
  buf x1155(s5892,s2091);
  buf x1156(s5900,s2085);
  buf x1157(s5908,s2335);
  buf x1158(s5916,s2329);
  buf x1159(s5924,s2323);
  nor x1160(s5969,s2091,s3731);
  buf x1161(s5988,s2111);
  buf x1162(s5996,s2105);
  buf x1163(s6004,s2099);
  buf x1164(s6012,s2085);
  buf x1165(s6020,s2335);
  buf x1166(s6028,s2329);
  buf x1167(s6036,s2323);
  buf x1168(s6044,s2091);
  nor x1169(s6057,s3731,s2091);
  buf x1170(s6439,s4175);
  buf x1171(s6447,s4172);
  buf x1172(s6455,s4169);
  buf x1173(s6463,s4163);
  buf x1174(s6471,s4160);
  buf x1175(s6474,s2175);
  buf x1176(s6479,s4157);
  buf x1177(s6482,s2171);
  buf x1178(s6487,s4154);
  buf x1179(s6490,s2167);
  buf x1180(s6495,s4166);
  buf x1181(s6503,s4151);
  buf x1182(s6506,s2163);
  buf x1183(s6570,s3838);
  buf x1184(s6578,s3833);
  buf x1185(s6586,s3828);
  buf x1186(s6594,s3821);
  buf x1187(s6602,s3816);
  buf x1188(s6610,s2198);
  buf x1189(s6618,s2192);
  buf x1190(s6626,s2186);
  buf x1191(s6634,s2179);
  nor x1192(s6671,s3821,s4422);
  buf x1193(s6721,s2179);
  buf x1194(s6729,s2192);
  buf x1195(s6732,s2186);
  buf x1196(s6737,s3816);
  buf x1197(s6740,s2198);
  buf x1198(s6745,s3828);
  buf x1199(s6748,s3821);
  buf x1200(s6755,s3838);
  buf x1201(s6758,s3833);
  buf x1202(s6765,s2320);
  buf x1203(s6773,s2329);
  buf x1204(s6776,s2323);
  buf x1205(s6781,s2085);
  buf x1206(s6784,s2335);
  buf x1207(s6789,s2099);
  buf x1208(s6792,s2091);
  buf x1209(s6799,s2111);
  buf x1210(s6802,s2105);
  nand x1211(s6832,s6719,s6720);
  buf x1212(s6856,s3838);
  buf x1213(s6864,s3833);
  buf x1214(s6872,s3828);
  buf x1215(s6880,s3816);
  buf x1216(s6888,s2198);
  buf x1217(s6896,s2192);
  buf x1218(s6904,s2186);
  buf x1219(s6912,s3821);
  buf x1220(s6920,s2179);
  nor x1221(s6925,s4422,s3821);
  nor x1222(s7041,s4396,s2179);
  buf x1223(s7205,s2163);
  buf x1224(s7213,s2171);
  buf x1225(s7216,s2167);
  buf x1226(s7224,s2175);
  not x1227(s7235,s7229);
  not x1228(s7236,s7232);
  not x1229(s7245,s7239);
  not x1230(s7246,s7242);
  buf x1231(s7265,s2065);
  buf x1232(s7273,s2073);
  buf x1233(s7276,s2069);
  buf x1234(s7283,s2081);
  buf x1235(s7286,s2077);
  not x1236(s7323,s7317);
  not x1237(s7324,s7320);
  not x1238(s7333,s7327);
  not x1239(s7334,s7330);
  buf x1240(s7361,s4511);
  buf x1241(s7364,s2081);
  buf x1242(s7369,s4508);
  buf x1243(s7372,s2077);
  buf x1244(s7377,s4505);
  buf x1245(s7380,s2073);
  buf x1246(s7385,s4499);
  buf x1247(s7388,s2065);
  buf x1248(s7393,s4496);
  buf x1249(s7401,s4493);
  buf x1250(s7409,s4490);
  buf x1251(s7417,s4502);
  buf x1252(s7420,s2069);
  buf x1253(s7428,s3695);
  not x1254(s7493,s7487);
  not x1255(s7494,s7490);
  not x1256(s7503,s7497);
  not x1257(s7504,s7500);
  buf x1258(s7515,s4493);
  buf x1259(s7518,s4490);
  buf x1260(s7523,s4499);
  buf x1261(s7526,s4496);
  buf x1262(s7531,s4505);
  buf x1263(s7534,s4502);
  buf x1264(s7541,s4511);
  buf x1265(s7544,s4508);
  buf x1266(s7551,s4151);
  buf x1267(s7559,s4157);
  buf x1268(s7562,s4154);
  buf x1269(s7567,s4163);
  buf x1270(s7570,s4160);
  buf x1271(s7575,s4169);
  buf x1272(s7578,s4166);
  buf x1273(s7585,s4175);
  buf x1274(s7588,s4172);
  nand x1275(s1176,s1121,s1112);
  nand x1276(s957,s912,s906);
  nand x1277(s791,s4881,s4888);
  nand x1278(s804,s4889,s4896);
  nand x1279(s826,s4897,s4904);
  nand x1280(s852,s4905,s4912);
  nand x1281(s894,s4921,s4928);
  nand x1282(s1025,s5191,s5198);
  nand x1283(s1037,s5199,s5206);
  nand x1284(s1054,s5207,s5214);
  nand x1285(s1073,s5215,s5222);
  nand x1286(s1092,s5223,s5230);
  nand x1287(s1154,s1152,s1153);
  nand x1288(s1158,s1156,s1157);
  nand x1289(s1215,s5250,s5253);
  nand x1290(s1224,s5258,s5261);
  nand x1291(s1225,s5255,s5262);
  nand x1292(s1233,s5266,s5269);
  nand x1293(s1234,s5263,s5270);
  nand x1294(s1238,s5284,s5287);
  nand x1295(s1247,s5292,s5295);
  nand x1296(s1248,s5289,s5296);
  nand x1297(s1256,s5300,s5303);
  nand x1298(s1257,s5297,s5304);
  nand x1299(s1261,s5318,s5321);
  nand x1300(s1270,s5326,s5329);
  nand x1301(s1271,s5323,s5330);
  nand x1302(s1279,s5334,s5337);
  nand x1303(s1280,s5331,s5338);
  nand x1304(s1545,s5393,s5400);
  nand x1305(s1555,s5401,s5408);
  nand x1306(s1572,s5409,s5416);
  nand x1307(s1597,s5417,s5424);
  nand x1308(s1608,s5425,s5432);
  nand x1309(s1629,s5433,s5440);
  nand x1310(s1654,s5441,s5448);
  nand x1311(s1686,s5449,s5456);
  nand x1312(s1694,s5457,s5464);
  nand x1313(s1794,s5745,s5752);
  nand x1314(s1804,s5753,s5760);
  nand x1315(s1821,s5761,s5768);
  nand x1316(s1849,s5769,s5776);
  nand x1317(s1858,s5777,s5784);
  nand x1318(s1868,s5785,s5792);
  nand x1319(s1884,s5793,s5800);
  nand x1320(s1902,s5801,s5808);
  nand x1321(s1920,s5809,s5816);
  nand x1322(s2954,s6370,s6373);
  nand x1323(s2955,s6367,s6374);
  nand x1324(s2963,s6378,s6381);
  nand x1325(s2964,s6375,s6382);
  nand x1326(s2971,s6386,s6389);
  nand x1327(s2972,s6383,s6390);
  nand x1328(s2980,s6394,s6397);
  nand x1329(s2981,s6391,s6398);
  nand x1330(s2990,s6402,s6405);
  nand x1331(s2991,s6399,s6406);
  nand x1332(s2999,s6410,s6413);
  nand x1333(s3000,s6407,s6414);
  nand x1334(s3007,s6418,s6421);
  nand x1335(s3008,s6415,s6422);
  nand x1336(s3016,s6426,s6429);
  nand x1337(s3017,s6423,s6430);
  nand x1338(s3019,s6434,s6437);
  nand x1339(s3020,s6431,s6438);
  nand x1340(s3174,s6522,s6525);
  nand x1341(s3175,s6519,s6526);
  nand x1342(s3184,s6530,s6533);
  nand x1343(s3185,s6527,s6534);
  nand x1344(s3193,s6538,s6541);
  nand x1345(s3194,s6535,s6542);
  nand x1346(s3201,s6546,s6549);
  nand x1347(s3202,s6543,s6550);
  nand x1348(s3213,s6562,s6565);
  nand x1349(s3214,s6559,s6566);
  not x1350(s3227,s3223);
  nand x1351(s3502,s6690,s6693);
  nand x1352(s3511,s6698,s6701);
  nand x1353(s3512,s6695,s6702);
  nand x1354(s3520,s6706,s6709);
  nand x1355(s3521,s6703,s6710);
  nand x1356(s4201,s7252,s7255);
  nand x1357(s4210,s7260,s7263);
  nand x1358(s4211,s7257,s7264);
  nand x1359(s4224,s7296,s7299);
  nand x1360(s4233,s7304,s7307);
  nand x1361(s4234,s7301,s7308);
  nand x1362(s4242,s7312,s7315);
  nand x1363(s4243,s7309,s7316);
  nand x1364(s4529,s7466,s7469);
  nand x1365(s4538,s7474,s7477);
  nand x1366(s4539,s7471,s7478);
  nand x1367(s4547,s7482,s7485);
  nand x1368(s4548,s7479,s7486);
  nand x1369(s4552,s7510,s7513);
  nand x1370(s4553,s7507,s7514);
  not x1371(s4946,s4942);
  nand x1372(s5347,s5342,s5345);
  nand x1373(s5348,s5339,s5346);
  nand x1374(s5357,s5352,s5355);
  nand x1375(s5358,s5349,s5356);
  nand x1376(s7237,s7232,s7235);
  nand x1377(s7238,s7229,s7236);
  nand x1378(s7247,s7242,s7245);
  nand x1379(s7248,s7239,s7246);
  nand x1380(s7325,s7320,s7323);
  nand x1381(s7326,s7317,s7324);
  nand x1382(s7335,s7330,s7333);
  nand x1383(s7336,s7327,s7334);
  nand x1384(s7495,s7490,s7493);
  nand x1385(s7496,s7487,s7494);
  nand x1386(s7505,s7500,s7503);
  nand x1387(s7506,s7497,s7504);
  nand x1388(s3244,s3227,s3220);
  nand x1389(s792,s790,s791);
  nand x1390(s805,s803,s804);
  nand x1391(s827,s825,s826);
  nand x1392(s853,s851,s852);
  nand x1393(s895,s893,s894);
  nand x1394(s1026,s1024,s1025);
  nand x1395(s1038,s1036,s1037);
  nand x1396(s1055,s1053,s1054);
  nand x1397(s1074,s1072,s1073);
  nand x1398(s1093,s1091,s1092);
  not x1399(s1155,s1154);
  nand x1400(s1217,s1215,s1216);
  nand x1401(s1226,s1224,s1225);
  nand x1402(s1235,s1233,s1234);
  nand x1403(s1240,s1238,s1239);
  nand x1404(s1249,s1247,s1248);
  nand x1405(s1258,s1256,s1257);
  nand x1406(s1263,s1261,s1262);
  nand x1407(s1272,s1270,s1271);
  nand x1408(s1281,s1279,s1280);
  not x1409(s5376,s5372);
  not x1410(s5384,s5380);
  nand x1411(s1546,s1544,s1545);
  nand x1412(s1556,s1554,s1555);
  nand x1413(s1573,s1571,s1572);
  nand x1414(s1598,s1596,s1597);
  nand x1415(s1609,s1607,s1608);
  nand x1416(s1630,s1628,s1629);
  nand x1417(s1655,s1653,s1654);
  nand x1418(s1687,s1685,s1686);
  nand x1419(s1695,s1693,s1694);
  nand x1420(s1795,s1793,s1794);
  nand x1421(s1805,s1803,s1804);
  nand x1422(s1822,s1820,s1821);
  nand x1423(s1850,s1848,s1849);
  nand x1424(s1859,s1857,s1858);
  nand x1425(s1869,s1867,s1868);
  nand x1426(s1885,s1883,s1884);
  nand x1427(s1903,s1901,s1902);
  nand x1428(s1921,s1919,s1920);
  not x1429(s5863,s5857);
  nand x1430(s2341,s5868,s5871);
  not x1431(s5872,s5868);
  nand x1432(s2352,s5876,s5879);
  not x1433(s5880,s5876);
  nand x1434(s2370,s5884,s5887);
  not x1435(s5888,s5884);
  nand x1436(s2398,s5892,s5895);
  not x1437(s5896,s5892);
  nand x1438(s2407,s5900,s5903);
  not x1439(s5904,s5900);
  nand x1440(s2418,s5908,s5911);
  not x1441(s5912,s5908);
  nand x1442(s2434,s5916,s5919);
  not x1443(s5920,s5916);
  nand x1444(s2452,s5924,s5927);
  not x1445(s5928,s5924);
  and x1446(s2481,s3682,s4389);
  not x1447(s5975,s5969);
  nand x1448(s2587,s5988,s5991);
  not x1449(s5992,s5988);
  nand x1450(s2598,s5996,s5999);
  not x1451(s6000,s5996);
  nand x1452(s2616,s6004,s6007);
  not x1453(s6008,s6004);
  nand x1454(s2641,s6012,s6015);
  not x1455(s6016,s6012);
  nand x1456(s2653,s6020,s6023);
  not x1457(s6024,s6020);
  nand x1458(s2674,s6028,s6031);
  not x1459(s6032,s6028);
  nand x1460(s2699,s6036,s6039);
  not x1461(s6040,s6036);
  and x1462(s2724,s3682,s4389);
  nand x1463(s2732,s6044,s6047);
  not x1464(s6048,s6044);
  nand x1465(s2956,s2954,s2955);
  nand x1466(s2965,s2963,s2964);
  nand x1467(s2973,s2971,s2972);
  nand x1468(s2982,s2980,s2981);
  nand x1469(s2992,s2990,s2991);
  nand x1470(s3001,s2999,s3000);
  nand x1471(s3009,s3007,s3008);
  nand x1472(s3018,s3016,s3017);
  nand x1473(s3021,s3019,s3020);
  not x1474(s6445,s6439);
  nand x1475(s3051,s6439,s6446);
  not x1476(s6453,s6447);
  nand x1477(s3061,s6447,s6454);
  not x1478(s6461,s6455);
  nand x1479(s3070,s6455,s6462);
  not x1480(s6469,s6463);
  nand x1481(s3081,s6463,s6470);
  not x1482(s6477,s6471);
  not x1483(s6478,s6474);
  not x1484(s6485,s6479);
  not x1485(s6486,s6482);
  not x1486(s6493,s6487);
  not x1487(s6494,s6490);
  not x1488(s6501,s6495);
  nand x1489(s3118,s6495,s6502);
  not x1490(s6509,s6503);
  not x1491(s6510,s6506);
  nand x1492(s3176,s3174,s3175);
  nand x1493(s3186,s3184,s3185);
  nand x1494(s3195,s3193,s3194);
  nand x1495(s3203,s3201,s3202);
  nand x1496(s3215,s3213,s3214);
  nand x1497(s3281,s6570,s6573);
  not x1498(s6574,s6570);
  nand x1499(s3293,s6578,s6581);
  not x1500(s6582,s6578);
  nand x1501(s3312,s6586,s6589);
  not x1502(s6590,s6586);
  nand x1503(s3342,s6594,s6597);
  not x1504(s6598,s6594);
  nand x1505(s3351,s6602,s6605);
  not x1506(s6606,s6602);
  nand x1507(s3363,s6610,s6613);
  not x1508(s6614,s6610);
  nand x1509(s3379,s6618,s6621);
  not x1510(s6622,s6618);
  nand x1511(s3397,s6626,s6629);
  not x1512(s6630,s6626);
  nand x1513(s3415,s6634,s6637);
  not x1514(s6638,s6634);
  not x1515(s6677,s6671);
  nand x1516(s3504,s3502,s3503);
  nand x1517(s3513,s3511,s3512);
  nand x1518(s3522,s3520,s3521);
  not x1519(s6727,s6721);
  nand x1520(s3526,s6721,s6728);
  not x1521(s6735,s6729);
  not x1522(s6736,s6732);
  not x1523(s6743,s6737);
  not x1524(s6744,s6740);
  not x1525(s6771,s6765);
  nand x1526(s3549,s6765,s6772);
  not x1527(s6779,s6773);
  not x1528(s6780,s6776);
  not x1529(s6787,s6781);
  not x1530(s6788,s6784);
  not x1531(s6836,s6832);
  nand x1532(s3843,s6856,s6859);
  not x1533(s6860,s6856);
  nand x1534(s3854,s6864,s6867);
  not x1535(s6868,s6864);
  nand x1536(s3872,s6872,s6875);
  not x1537(s6876,s6872);
  nand x1538(s3897,s6880,s6883);
  not x1539(s6884,s6880);
  nand x1540(s3909,s6888,s6891);
  not x1541(s6892,s6888);
  nand x1542(s3930,s6896,s6899);
  not x1543(s6900,s6896);
  nand x1544(s3955,s6904,s6907);
  not x1545(s6908,s6904);
  nand x1546(s3987,s6912,s6915);
  not x1547(s6916,s6912);
  nand x1548(s3995,s6920,s6923);
  not x1549(s6924,s6920);
  not x1550(s7211,s7205);
  nand x1551(s4179,s7205,s7212);
  not x1552(s7219,s7213);
  not x1553(s7220,s7216);
  nand x1554(s4196,s7224,s7227);
  not x1555(s7228,s7224);
  nand x1556(s4203,s4201,s4202);
  nand x1557(s4212,s4210,s4211);
  not x1558(s7271,s7265);
  nand x1559(s4220,s7265,s7272);
  nand x1560(s4226,s4224,s4225);
  nand x1561(s4235,s4233,s4234);
  nand x1562(s4244,s4242,s4243);
  not x1563(s7367,s7361);
  not x1564(s7368,s7364);
  not x1565(s7375,s7369);
  not x1566(s7376,s7372);
  not x1567(s7383,s7377);
  not x1568(s7384,s7380);
  not x1569(s7391,s7385);
  not x1570(s7392,s7388);
  not x1571(s7399,s7393);
  nand x1572(s4326,s7393,s7400);
  not x1573(s7407,s7401);
  nand x1574(s4335,s7401,s7408);
  not x1575(s7415,s7409);
  nand x1576(s4343,s7409,s7416);
  not x1577(s7423,s7417);
  not x1578(s7424,s7420);
  nand x1579(s4353,s7428,s7431);
  not x1580(s7432,s7428);
  nand x1581(s4531,s4529,s4530);
  nand x1582(s4540,s4538,s4539);
  nand x1583(s4549,s4547,s4548);
  nand x1584(s4554,s4552,s4553);
  not x1585(s7521,s7515);
  not x1586(s7522,s7518);
  not x1587(s7529,s7523);
  not x1588(s7530,s7526);
  not x1589(s7557,s7551);
  nand x1590(s4576,s7551,s7558);
  not x1591(s7565,s7559);
  not x1592(s7566,s7562);
  not x1593(s7573,s7567);
  not x1594(s7574,s7570);
  not x1595(s4936,s4932);
  nand x1596(s4937,s4932,s4935);
  not x1597(s4977,s4973);
  nand x1598(s4978,s4973,s4976);
  not x1599(s5105,s5099);
  nand x1600(s5359,s5357,s5358);
  nand x1601(s5362,s5347,s5348);
  not x1602(s5529,s5523);
  not x1603(s5675,s5669);
  buf x1604(s5932,s4389);
  buf x1605(s5977,s2391);
  buf x1606(s6052,s4389);
  not x1607(s6063,s6057);
  buf x1608(s6115,s2635);
  nor x1609(s6173,s3682,s4389);
  buf x1610(s6679,s3335);
  not x1611(s6751,s6745);
  not x1612(s6752,s6748);
  not x1613(s6761,s6755);
  not x1614(s6762,s6758);
  not x1615(s6795,s6789);
  not x1616(s6796,s6792);
  not x1617(s6805,s6799);
  not x1618(s6806,s6802);
  not x1619(s6931,s6925);
  buf x1620(s6983,s3891);
  not x1621(s7047,s7041);
  buf x1622(s7129,s3979);
  not x1623(s7279,s7273);
  not x1624(s7280,s7276);
  not x1625(s7289,s7283);
  not x1626(s7290,s7286);
  nand x1627(s7337,s7247,s7248);
  nand x1628(s7340,s7237,s7238);
  nand x1629(s7353,s7335,s7336);
  nand x1630(s7356,s7325,s7326);
  not x1631(s7537,s7531);
  not x1632(s7538,s7534);
  not x1633(s7547,s7541);
  not x1634(s7548,s7544);
  not x1635(s7581,s7575);
  not x1636(s7582,s7578);
  not x1637(s7591,s7585);
  not x1638(s7592,s7588);
  nand x1639(s7595,s7505,s7506);
  nand x1640(s7598,s7495,s7496);
  nand x1641(s2342,s5865,s5872);
  nand x1642(s2353,s5873,s5880);
  nand x1643(s2371,s5881,s5888);
  nand x1644(s2399,s5889,s5896);
  nand x1645(s2408,s5897,s5904);
  nand x1646(s2419,s5905,s5912);
  nand x1647(s2435,s5913,s5920);
  nand x1648(s2453,s5921,s5928);
  nand x1649(s2588,s5985,s5992);
  nand x1650(s2599,s5993,s6000);
  nand x1651(s2617,s6001,s6008);
  nand x1652(s2642,s6009,s6016);
  nand x1653(s2654,s6017,s6024);
  nand x1654(s2675,s6025,s6032);
  nand x1655(s2700,s6033,s6040);
  nand x1656(s2733,s6041,s6048);
  nand x1657(s3050,s6442,s6445);
  nand x1658(s3060,s6450,s6453);
  nand x1659(s3069,s6458,s6461);
  nand x1660(s3080,s6466,s6469);
  nand x1661(s3091,s6474,s6477);
  nand x1662(s3092,s6471,s6478);
  nand x1663(s3100,s6482,s6485);
  nand x1664(s3101,s6479,s6486);
  nand x1665(s3108,s6490,s6493);
  nand x1666(s3109,s6487,s6494);
  nand x1667(s3117,s6498,s6501);
  nand x1668(s3120,s6506,s6509);
  nand x1669(s3121,s6503,s6510);
  nand x1670(s3282,s6567,s6574);
  nand x1671(s3294,s6575,s6582);
  nand x1672(s3313,s6583,s6590);
  nand x1673(s3343,s6591,s6598);
  nand x1674(s3352,s6599,s6606);
  nand x1675(s3364,s6607,s6614);
  nand x1676(s3380,s6615,s6622);
  nand x1677(s3398,s6623,s6630);
  nand x1678(s3416,s6631,s6638);
  nand x1679(s3525,s6724,s6727);
  nand x1680(s3534,s6732,s6735);
  nand x1681(s3535,s6729,s6736);
  nand x1682(s3543,s6740,s6743);
  nand x1683(s3544,s6737,s6744);
  nand x1684(s3548,s6768,s6771);
  nand x1685(s3557,s6776,s6779);
  nand x1686(s3558,s6773,s6780);
  nand x1687(s3566,s6784,s6787);
  nand x1688(s3567,s6781,s6788);
  nand x1689(s3844,s6853,s6860);
  nand x1690(s3855,s6861,s6868);
  nand x1691(s3873,s6869,s6876);
  nand x1692(s3898,s6877,s6884);
  nand x1693(s3910,s6885,s6892);
  nand x1694(s3931,s6893,s6900);
  nand x1695(s3956,s6901,s6908);
  nand x1696(s3988,s6909,s6916);
  nand x1697(s3996,s6917,s6924);
  nand x1698(s4178,s7208,s7211);
  nand x1699(s4187,s7216,s7219);
  nand x1700(s4188,s7213,s7220);
  nand x1701(s4197,s7221,s7228);
  nand x1702(s4219,s7268,s7271);
  nand x1703(s4289,s7364,s7367);
  nand x1704(s4290,s7361,s7368);
  nand x1705(s4298,s7372,s7375);
  nand x1706(s4299,s7369,s7376);
  nand x1707(s4306,s7380,s7383);
  nand x1708(s4307,s7377,s7384);
  nand x1709(s4315,s7388,s7391);
  nand x1710(s4316,s7385,s7392);
  nand x1711(s4325,s7396,s7399);
  nand x1712(s4334,s7404,s7407);
  nand x1713(s4342,s7412,s7415);
  nand x1714(s4350,s7420,s7423);
  nand x1715(s4351,s7417,s7424);
  nand x1716(s4354,s7425,s7432);
  nand x1717(s4561,s7518,s7521);
  nand x1718(s4562,s7515,s7522);
  nand x1719(s4570,s7526,s7529);
  nand x1720(s4571,s7523,s7530);
  nand x1721(s4575,s7554,s7557);
  nand x1722(s4584,s7562,s7565);
  nand x1723(s4585,s7559,s7566);
  nand x1724(s4593,s7570,s7573);
  nand x1725(s4594,s7567,s7574);
  nand x1726(s4938,s4929,s4936);
  nand x1727(s4979,s4970,s4977);
  nand x1728(s6753,s6748,s6751);
  nand x1729(s6754,s6745,s6752);
  nand x1730(s6763,s6758,s6761);
  nand x1731(s6764,s6755,s6762);
  nand x1732(s6797,s6792,s6795);
  nand x1733(s6798,s6789,s6796);
  nand x1734(s6807,s6802,s6805);
  nand x1735(s6808,s6799,s6806);
  nand x1736(s7281,s7276,s7279);
  nand x1737(s7282,s7273,s7280);
  nand x1738(s7291,s7286,s7289);
  nand x1739(s7292,s7283,s7290);
  nand x1740(s7539,s7534,s7537);
  nand x1741(s7540,s7531,s7538);
  nand x1742(s7549,s7544,s7547);
  nand x1743(s7550,s7541,s7548);
  nand x1744(s7583,s7578,s7581);
  nand x1745(s7584,s7575,s7582);
  nand x1746(s7593,s7588,s7591);
  nand x1747(s7594,s7585,s7592);
  not x1748(s1856,s1850);
  and x1749(s920,s895,s853,s827,s805,s792);
  and x1750(s925,s792,s821);
  and x1751(s926,s805,s792,s845);
  and x1752(s927,s827,s792,s868,s805);
  and x1753(s928,s853,s827,s792,s877,s805);
  and x1754(s937,s805,s845);
  and x1755(s938,s827,s868,s805);
  and x1756(s939,s853,s827,s877,s805);
  and x1757(s940,s895,s827,s805,s853);
  and x1758(s941,s805,s845);
  and x1759(s942,s827,s868,s805);
  and x1760(s943,s853,s827,s877,s805);
  and x1761(s944,s827,s868);
  and x1762(s945,s853,s827,s877);
  and x1763(s946,s895,s827,s853);
  and x1764(s947,s827,s868);
  and x1765(s948,s853,s827,s877);
  and x1766(s949,s853,s877);
  and x1767(s956,s895,s853);
  and x1768(s1122,s1038,s1093,s1055,s1026,s1074);
  and x1769(s1125,s1026,s1050);
  and x1770(s1126,s1038,s1026,s1068);
  and x1771(s1127,s1055,s1026,s1086,s1038);
  and x1772(s1128,s1074,s1055,s1026,s1102,s1038);
  and x1773(s1132,s1038,s1068);
  and x1774(s1133,s1055,s1086,s1038);
  and x1775(s1134,s1074,s1055,s1102,s1038);
  and x1776(s1137,s1086,s1055);
  and x1777(s1138,s1074,s1055,s1102);
  and x1778(s1141,s1074,s1102);
  not x1779(s1221,s1217);
  not x1780(s1230,s1226);
  not x1781(s1244,s1240);
  not x1782(s1253,s1249);
  not x1783(s1267,s1263);
  not x1784(s1276,s1272);
  buf x1785(s1284,s1235);
  buf x1786(s1288,s1235);
  buf x1787(s1292,s1258);
  buf x1788(s1296,s1258);
  buf x1789(s1300,s1281);
  buf x1790(s1304,s1281);
  and x1791(s1702,s1687,s1573,s1556,s1546);
  and x1792(s1705,s1546,s1567);
  and x1793(s1706,s1556,s1546,s1584);
  and x1794(s1707,s1573,s1546,s1590,s1556);
  and x1795(s1709,s1556,s1584);
  and x1796(s1710,s1573,s1590,s1556);
  and x1797(s1711,s1687,s1573,s1556);
  and x1798(s1712,s1556,s1584);
  and x1799(s1713,s1573,s1590,s1556);
  and x1800(s1714,s1573,s1590);
  and x1801(s1718,s1695,s1655,s1630,s1609,s1598);
  and x1802(s1722,s1598,s1624);
  and x1803(s1723,s1609,s1598,s1647);
  and x1804(s1724,s1630,s1598,s1669,s1609);
  and x1805(s1725,s1655,s1630,s1598,s1677,s1609);
  and x1806(s1733,s1609,s1647);
  and x1807(s1734,s1630,s1669,s1609);
  and x1808(s1735,s1655,s1630,s1677,s1609);
  and x1809(s1736,s1695,s1630,s1609,s1655);
  and x1810(s1737,s1609,s1647);
  and x1811(s1738,s1630,s1669,s1609);
  and x1812(s1739,s1655,s1630,s1677,s1609);
  and x1813(s1740,s1630,s1669);
  and x1814(s1741,s1655,s1630,s1677);
  and x1815(s1742,s1695,s1630,s1655);
  and x1816(s1743,s1630,s1669);
  and x1817(s1744,s1655,s1630,s1677);
  and x1818(s1745,s1655,s1677);
  and x1819(s1749,s1687,s1573);
  and x1820(s1750,s1695,s1655);
  and x1821(s1935,s1805,s1850,s1822,s1795);
  and x1822(s1938,s1795,s1816);
  and x1823(s1939,s1805,s1795,s1834);
  and x1824(s1940,s1822,s1795,s1841,s1805);
  and x1825(s1942,s1805,s1834);
  and x1826(s1943,s1822,s1841,s1805);
  and x1827(s1944,s1850,s1822,s1805);
  and x1828(s1945,s1805,s1834);
  and x1829(s1946,s1841,s1822,s1805);
  and x1830(s1947,s1822,s1841);
  and x1831(s1948,s1850,s1822);
  and x1832(s1949,s1822,s1841);
  and x1833(s1950,s1869,s1921,s1885,s1859,s1903);
  and x1834(s1953,s1859,s1880);
  and x1835(s1954,s1869,s1859,s1897);
  and x1836(s1955,s1885,s1859,s1914,s1869);
  and x1837(s1956,s1903,s1885,s1859,s1929,s1869);
  and x1838(s1960,s1869,s1897);
  and x1839(s1961,s1885,s1914,s1869);
  and x1840(s1962,s1903,s1885,s1929,s1869);
  and x1841(s1965,s1914,s1885);
  and x1842(s1966,s1903,s1885,s1929);
  and x1843(s1969,s1903,s1929);
  nand x1844(s2343,s2341,s2342);
  nand x1845(s2354,s2352,s2353);
  nand x1846(s2372,s2370,s2371);
  nand x1847(s2400,s2398,s2399);
  nand x1848(s2409,s2407,s2408);
  nand x1849(s2420,s2418,s2419);
  nand x1850(s2436,s2434,s2435);
  nand x1851(s2454,s2452,s2453);
  nand x1852(s2470,s5932,s5935);
  not x1853(s5936,s5932);
  not x1854(s5983,s5977);
  nand x1855(s2589,s2587,s2588);
  nand x1856(s2600,s2598,s2599);
  nand x1857(s2618,s2616,s2617);
  nand x1858(s2643,s2641,s2642);
  nand x1859(s2655,s2653,s2654);
  nand x1860(s2676,s2674,s2675);
  nand x1861(s2701,s2699,s2700);
  nand x1862(s2734,s2732,s2733);
  nand x1863(s2740,s6052,s6055);
  not x1864(s6056,s6052);
  and x1865(s3022,s3018,s2973,s2965,s2956);
  and x1866(s3025,s2956,s2970);
  and x1867(s3026,s2965,s2956,s2977);
  and x1868(s3027,s2973,s2956,s2979,s2965);
  and x1869(s3029,s3021,s3009,s3001,s2992,s2982);
  and x1870(s3030,s2982,s2998);
  and x1871(s3031,s2992,s2982,s3006);
  and x1872(s3032,s3001,s2982,s3013,s2992);
  and x1873(s3033,s3009,s3001,s2982,s3015,s2992);
  nand x1874(s3052,s3050,s3051);
  nand x1875(s3062,s3060,s3061);
  nand x1876(s3071,s3069,s3070);
  nand x1877(s3082,s3080,s3081);
  nand x1878(s3093,s3091,s3092);
  nand x1879(s3102,s3100,s3101);
  nand x1880(s3110,s3108,s3109);
  nand x1881(s3119,s3117,s3118);
  nand x1882(s3122,s3120,s3121);
  and x1883(s3228,s3215,s3203,s3195,s3186,s3176);
  and x1884(s3231,s3176,s3192);
  and x1885(s3232,s3186,s3176,s3200);
  and x1886(s3233,s3195,s3176,s3207,s3186);
  and x1887(s3234,s3203,s3195,s3176,s3209,s3186);
  nand x1888(s3283,s3281,s3282);
  nand x1889(s3295,s3293,s3294);
  nand x1890(s3314,s3312,s3313);
  nand x1891(s3344,s3342,s3343);
  nand x1892(s3353,s3351,s3352);
  nand x1893(s3365,s3363,s3364);
  nand x1894(s3381,s3379,s3380);
  nand x1895(s3399,s3397,s3398);
  nand x1896(s3417,s3415,s3416);
  not x1897(s6685,s6679);
  not x1898(s3508,s3504);
  not x1899(s3517,s3513);
  nand x1900(s3527,s3525,s3526);
  nand x1901(s3536,s3534,s3535);
  nand x1902(s3545,s3543,s3544);
  nand x1903(s3550,s3548,s3549);
  nand x1904(s3559,s3557,s3558);
  nand x1905(s3568,s3566,s3567);
  buf x1906(s3571,s3522);
  buf x1907(s3575,s3522);
  nand x1908(s3845,s3843,s3844);
  nand x1909(s3856,s3854,s3855);
  nand x1910(s3874,s3872,s3873);
  nand x1911(s3899,s3897,s3898);
  nand x1912(s3911,s3909,s3910);
  nand x1913(s3932,s3930,s3931);
  nand x1914(s3957,s3955,s3956);
  nand x1915(s3989,s3987,s3988);
  nand x1916(s3997,s3995,s3996);
  nand x1917(s4180,s4178,s4179);
  nand x1918(s4189,s4187,s4188);
  nand x1919(s4198,s4196,s4197);
  not x1920(s4207,s4203);
  not x1921(s4216,s4212);
  nand x1922(s4221,s4219,s4220);
  not x1923(s4230,s4226);
  not x1924(s4239,s4235);
  buf x1925(s4263,s4244);
  buf x1926(s4267,s4244);
  nand x1927(s4291,s4289,s4290);
  nand x1928(s4300,s4298,s4299);
  nand x1929(s4308,s4306,s4307);
  nand x1930(s4317,s4315,s4316);
  nand x1931(s4327,s4325,s4326);
  nand x1932(s4336,s4334,s4335);
  nand x1933(s4344,s4342,s4343);
  nand x1934(s4352,s4350,s4351);
  nand x1935(s4355,s4353,s4354);
  not x1936(s4535,s4531);
  not x1937(s4544,s4540);
  not x1938(s4558,s4554);
  nand x1939(s4563,s4561,s4562);
  nand x1940(s4572,s4570,s4571);
  nand x1941(s4577,s4575,s4576);
  nand x1942(s4586,s4584,s4585);
  nand x1943(s4595,s4593,s4594);
  buf x1944(s4598,s4549);
  buf x1945(s4602,s4549);
  buf x1946(s4716,s1921);
  buf x1947(s4724,s1859);
  buf x1948(s4732,s1869);
  buf x1949(s4740,s1885);
  buf x1950(s4748,s1903);
  buf x1951(s4756,s1093);
  buf x1952(s4764,s1026);
  buf x1953(s4772,s1038);
  buf x1954(s4780,s1055);
  buf x1955(s4788,s1074);
  nand x1956(s4939,s4937,s4938);
  nand x1957(s4980,s4978,s4979);
  buf x1958(s5044,s895);
  buf x1959(s5054,s853);
  buf x1960(s5064,s792);
  buf x1961(s5074,s827);
  buf x1962(s5084,s805);
  buf x1963(s5094,s805);
  buf x1964(s5132,s895);
  buf x1965(s5142,s853);
  buf x1966(s5152,s792);
  buf x1967(s5162,s827);
  not x1968(s5365,s5359);
  not x1969(s5366,s5362);
  buf x1970(s5488,s1687);
  buf x1971(s5498,s1573);
  buf x1972(s5508,s1546);
  buf x1973(s5518,s1556);
  buf x1974(s5546,s1687);
  buf x1975(s5556,s1573);
  buf x1976(s5566,s1546);
  buf x1977(s5576,s1556);
  buf x1978(s5614,s1695);
  buf x1979(s5624,s1655);
  buf x1980(s5634,s1598);
  buf x1981(s5644,s1630);
  buf x1982(s5654,s1609);
  buf x1983(s5664,s1609);
  buf x1984(s5702,s1695);
  buf x1985(s5712,s1655);
  buf x1986(s5722,s1598);
  buf x1987(s5732,s1630);
  buf x1988(s5820,s1795);
  buf x1989(s5828,s1795);
  buf x1990(s5836,s1805);
  buf x1991(s5844,s1805);
  buf x1992(s5852,s1822);
  buf x1993(s5860,s1822);
  not x1994(s6121,s6115);
  not x1995(s6179,s6173);
  buf x1996(s6261,s2724);
  not x1997(s7359,s7353);
  not x1998(s7360,s7356);
  not x1999(s7343,s7337);
  not x2000(s7344,s7340);
  nand x2001(s6809,s6763,s6764);
  nand x2002(s6812,s6753,s6754);
  nand x2003(s6819,s6807,s6808);
  nand x2004(s6822,s6797,s6798);
  not x2005(s6989,s6983);
  not x2006(s7135,s7129);
  nand x2007(s7345,s7291,s7292);
  nand x2008(s7348,s7281,s7282);
  not x2009(s7601,s7595);
  not x2010(s7602,s7598);
  nand x2011(s7603,s7549,s7550);
  nand x2012(s7606,s7539,s7540);
  nand x2013(s7611,s7593,s7594);
  nand x2014(s7614,s7583,s7584);
  or x2015(s929,s802,s925,s926,s927,s928);
  or x2016(s950,s868,s949);
  or x2017(s1129,s1035,s1125,s1126,s1127,s1128);
  or x2018(s1708,s1553,s1705,s1706,s1707);
  or x2019(s1715,s1584,s1714);
  or x2020(s1726,s1606,s1722,s1723,s1724,s1725);
  or x2021(s1746,s1669,s1745);
  or x2022(s1941,s1802,s1938,s1939,s1940);
  or x2023(s1957,s1866,s1953,s1954,s1955,s1956);
  nand x2024(s2471,s5929,s5936);
  nand x2025(s2741,s6049,s6056);
  or x2026(s3028,s2962,s3025,s3026,s3027);
  or x2027(s3034,s2989,s3030,s3031,s3032,s3033);
  or x2028(s3235,s3183,s3231,s3232,s3233,s3234);
  or x2029(s5014,s845,s944,s945,s946);
  or x2030(s5034,s821,s937,s938,s939,s940);
  nor x2031(s5102,s845,s947,s948);
  nor x2032(s5122,s821,s941,s942,s943);
  nand x2033(s5367,s5362,s5365);
  nand x2034(s5368,s5359,s5366);
  or x2035(s5478,s1567,s1709,s1710,s1711);
  nor x2036(s5536,s1567,s1712,s1713);
  or x2037(s5584,s1647,s1740,s1741,s1742);
  or x2038(s5604,s1624,s1733,s1734,s1735,s1736);
  nor x2039(s5672,s1647,s1743,s1744);
  nor x2040(s5692,s1624,s1737,s1738,s1739);
  or x2041(s5817,s1816,s1942,s1943,s1944);
  nor x2042(s5825,s1816,s1945,s1946);
  or x2043(s5833,s1834,s1947,s1948);
  nor x2044(s5841,s1834,s1949);
  nand x2045(s6340,s7356,s7359);
  nand x2046(s6341,s7353,s7360);
  nand x2047(s6350,s7340,s7343);
  nand x2048(s6351,s7337,s7344);
  nand x2049(s7436,s7598,s7601);
  nand x2050(s7437,s7595,s7602);
  not x2051(s4720,s4716);
  not x2052(s4728,s4724);
  not x2053(s4736,s4732);
  not x2054(s4744,s4740);
  not x2055(s4752,s4748);
  not x2056(s4760,s4756);
  not x2057(s4768,s4764);
  not x2058(s4776,s4772);
  not x2059(s4784,s4780);
  not x2060(s4792,s4788);
  not x2061(s3350,s3344);
  not x2062(s2406,s2400);
  not x2063(s924,s920);
  not x2064(s5088,s5084);
  not x2065(s5098,s5094);
  and x2066(s997,s902,s920);
  and x2067(s1146,s1108,s1122);
  not x2068(s1287,s1284);
  not x2069(s1291,s1288);
  not x2070(s1295,s1292);
  not x2071(s1299,s1296);
  not x2072(s1303,s1300);
  not x2073(s1307,s1304);
  and x2074(s1309,s1226,s1217,s1284);
  and x2075(s1312,s1230,s1221,s1288);
  and x2076(s1315,s1249,s1240,s1292);
  and x2077(s1318,s1253,s1244,s1296);
  and x2078(s1321,s1272,s1263,s1300);
  and x2079(s1324,s1276,s1267,s1304);
  not x2080(s1721,s1718);
  not x2081(s5522,s5518);
  not x2082(s5580,s5576);
  not x2083(s5658,s5654);
  not x2084(s5668,s5664);
  and x2085(s1788,s1702,s1718);
  and x2086(s1974,s1935,s1950);
  not x2087(s5824,s5820);
  not x2088(s5832,s5828);
  not x2089(s5840,s5836);
  not x2090(s5848,s5844);
  nand x2091(s1999,s5852,s5855);
  not x2092(s5856,s5852);
  nand x2093(s2003,s5860,s5863);
  not x2094(s5864,s5860);
  nand x2095(s2472,s2470,s2471);
  and x2096(s2487,s2354,s2400,s2372,s2343);
  and x2097(s2492,s2343,s2366);
  and x2098(s2493,s2354,s2343,s2384);
  and x2099(s2494,s2372,s2343,s2391,s2354);
  and x2100(s2500,s2354,s2384);
  and x2101(s2501,s2372,s2391,s2354);
  and x2102(s2502,s2400,s2372,s2354);
  and x2103(s2503,s2354,s2384);
  and x2104(s2504,s2391,s2372,s2354);
  and x2105(s2505,s2372,s2391);
  and x2106(s2506,s2400,s2372);
  and x2107(s2507,s2372,s2391);
  and x2108(s2511,s2409,s2431);
  and x2109(s2512,s2420,s2409,s2448);
  and x2110(s2513,s2436,s2409,s2465,s2420);
  and x2111(s2514,s2454,s2436,s2409,s2481,s2420);
  and x2112(s2518,s2420,s2448);
  and x2113(s2519,s2436,s2465,s2420);
  and x2114(s2520,s2454,s2436,s2481,s2420);
  and x2115(s2523,s2465,s2436);
  and x2116(s2524,s2454,s2436,s2481);
  and x2117(s2527,s2454,s2481);
  nand x2118(s2742,s2740,s2741);
  and x2119(s2749,s2734,s2618,s2600,s2589);
  and x2120(s2754,s2589,s2612);
  and x2121(s2755,s2600,s2589,s2629);
  and x2122(s2756,s2618,s2589,s2635,s2600);
  and x2123(s2762,s2600,s2629);
  and x2124(s2763,s2618,s2635,s2600);
  and x2125(s2764,s2734,s2618,s2600);
  and x2126(s2765,s2600,s2629);
  and x2127(s2766,s2618,s2635,s2600);
  and x2128(s2767,s2618,s2635);
  and x2129(s2776,s2643,s2670);
  and x2130(s2777,s2655,s2643,s2693);
  and x2131(s2778,s2676,s2643,s2715,s2655);
  and x2132(s2779,s2701,s2676,s2643,s2724,s2655);
  and x2133(s2788,s2655,s2693);
  and x2134(s2789,s2676,s2715,s2655);
  and x2135(s2790,s2701,s2676,s2724,s2655);
  and x2136(s2792,s2655,s2693);
  and x2137(s2793,s2676,s2715,s2655);
  and x2138(s2794,s2701,s2676,s2724,s2655);
  and x2139(s2795,s2676,s2715);
  and x2140(s2796,s2701,s2676,s2724);
  and x2141(s2798,s2676,s2715);
  and x2142(s2799,s2701,s2676,s2724);
  and x2143(s2800,s2701,s2724);
  and x2144(s2804,s2734,s2618);
  and x2145(s3035,s3022,s3029);
  and x2146(s3045,s3022,s3034);
  and x2147(s3123,s3119,s3071,s3062,s3052);
  and x2148(s3128,s3052,s3068);
  and x2149(s3129,s3062,s3052,s3076);
  and x2150(s3130,s3071,s3052,s3079,s3062);
  and x2151(s3136,s3122,s3110,s3102,s3093,s3082);
  and x2152(s3139,s3082,s3099);
  and x2153(s3140,s3093,s3082,s3107);
  and x2154(s3141,s3102,s3082,s3114,s3093);
  and x2155(s3142,s3110,s3102,s3082,s3116,s3093);
  and x2156(s3249,s3216,s3228);
  and x2157(s3431,s3295,s3344,s3314,s3283);
  and x2158(s3434,s3283,s3308);
  and x2159(s3435,s3295,s3283,s3327);
  and x2160(s3436,s3314,s3283,s3335,s3295);
  and x2161(s3438,s3295,s3327);
  and x2162(s3439,s3314,s3335,s3295);
  and x2163(s3440,s3344,s3314,s3295);
  and x2164(s3441,s3295,s3327);
  and x2165(s3442,s3335,s3314,s3295);
  and x2166(s3443,s3314,s3335);
  and x2167(s3444,s3344,s3314);
  and x2168(s3445,s3314,s3335);
  and x2169(s3446,s3365,s3417,s3381,s3353,s3399);
  and x2170(s3449,s3353,s3376);
  and x2171(s3450,s3365,s3353,s3393);
  and x2172(s3451,s3381,s3353,s3410,s3365);
  and x2173(s3452,s3399,s3381,s3353,s3425,s3365);
  and x2174(s3456,s3365,s3393);
  and x2175(s3457,s3381,s3410,s3365);
  and x2176(s3458,s3399,s3381,s3425,s3365);
  and x2177(s3460,s3410,s3381);
  and x2178(s3461,s3399,s3381,s3425);
  and x2179(s3463,s3399,s3425);
  not x2180(s3531,s3527);
  not x2181(s3540,s3536);
  not x2182(s3554,s3550);
  not x2183(s3563,s3559);
  not x2184(s3574,s3571);
  not x2185(s3578,s3575);
  buf x2186(s3579,s3545);
  buf x2187(s3583,s3545);
  buf x2188(s3587,s3568);
  buf x2189(s3591,s3568);
  and x2190(s3596,s3513,s3504,s3571);
  and x2191(s3599,s3517,s3508,s3575);
  and x2192(s4004,s3989,s3874,s3856,s3845);
  and x2193(s4007,s3845,s3868);
  and x2194(s4008,s3856,s3845,s3885);
  and x2195(s4009,s3874,s3845,s3891,s3856);
  and x2196(s4011,s3856,s3885);
  and x2197(s4012,s3874,s3891,s3856);
  and x2198(s4013,s3989,s3874,s3856);
  and x2199(s4014,s3856,s3885);
  and x2200(s4015,s3874,s3891,s3856);
  and x2201(s4016,s3874,s3891);
  and x2202(s4020,s3997,s3957,s3932,s3911,s3899);
  and x2203(s4024,s3899,s3926);
  and x2204(s4025,s3911,s3899,s3949);
  and x2205(s4026,s3932,s3899,s3971,s3911);
  and x2206(s4027,s3957,s3932,s3899,s3979,s3911);
  and x2207(s4035,s3911,s3949);
  and x2208(s4036,s3932,s3971,s3911);
  and x2209(s4037,s3957,s3932,s3979,s3911);
  and x2210(s4038,s3997,s3932,s3911,s3957);
  and x2211(s4039,s3911,s3949);
  and x2212(s4040,s3932,s3971,s3911);
  and x2213(s4041,s3957,s3932,s3979,s3911);
  and x2214(s4042,s3932,s3971);
  and x2215(s4043,s3957,s3932,s3979);
  and x2216(s4044,s3997,s3932,s3957);
  and x2217(s4045,s3932,s3971);
  and x2218(s4046,s3957,s3932,s3979);
  and x2219(s4047,s3957,s3979);
  and x2220(s4051,s3989,s3874);
  and x2221(s4052,s3997,s3957);
  not x2222(s4184,s4180);
  not x2223(s4193,s4189);
  buf x2224(s4247,s4198);
  buf x2225(s4251,s4198);
  buf x2226(s4255,s4221);
  buf x2227(s4259,s4221);
  not x2228(s4266,s4263);
  not x2229(s4270,s4267);
  and x2230(s4284,s4235,s4226,s4263);
  and x2231(s4287,s4239,s4230,s4267);
  and x2232(s4356,s4352,s4308,s4300,s4291);
  and x2233(s4361,s4291,s4305);
  and x2234(s4362,s4300,s4291,s4312);
  and x2235(s4363,s4308,s4291,s4314,s4300);
  and x2236(s4369,s4355,s4344,s4336,s4327,s4317);
  and x2237(s4372,s4317,s4333);
  and x2238(s4373,s4327,s4317,s4341);
  and x2239(s4374,s4336,s4317,s4348,s4327);
  and x2240(s4375,s4344,s4336,s4317,s4349,s4327);
  not x2241(s4567,s4563);
  not x2242(s4581,s4577);
  not x2243(s4590,s4586);
  not x2244(s4601,s4598);
  not x2245(s4605,s4602);
  buf x2246(s4606,s4572);
  buf x2247(s4610,s4572);
  buf x2248(s4614,s4595);
  buf x2249(s4618,s4595);
  and x2250(s4623,s4540,s4531,s4598);
  and x2251(s4626,s4544,s4535,s4602);
  buf x2252(s4796,s3417);
  buf x2253(s4804,s3353);
  buf x2254(s4812,s3365);
  buf x2255(s4820,s3381);
  buf x2256(s4828,s3399);
  buf x2257(s4844,s2409);
  buf x2258(s4852,s2420);
  buf x2259(s4860,s2436);
  buf x2260(s4868,s2454);
  not x2261(s4945,s4939);
  nand x2262(s4948,s4939,s4946);
  not x2263(s4986,s4980);
  nand x2264(s4989,s4980,s4987);
  not x2265(s5048,s5044);
  not x2266(s5058,s5054);
  not x2267(s5068,s5064);
  not x2268(s5078,s5074);
  not x2269(s5166,s5162);
  not x2270(s5136,s5132);
  not x2271(s5146,s5142);
  not x2272(s5156,s5152);
  nand x2273(s5388,s5367,s5368);
  not x2274(s5492,s5488);
  not x2275(s5502,s5498);
  not x2276(s5512,s5508);
  not x2277(s5550,s5546);
  not x2278(s5560,s5556);
  not x2279(s5570,s5566);
  not x2280(s5618,s5614);
  not x2281(s5628,s5624);
  not x2282(s5638,s5634);
  not x2283(s5648,s5644);
  not x2284(s5736,s5732);
  not x2285(s5706,s5702);
  not x2286(s5716,s5712);
  not x2287(s5726,s5722);
  buf x2288(s5940,s2343);
  buf x2289(s5948,s2343);
  buf x2290(s5956,s2354);
  buf x2291(s5964,s2354);
  buf x2292(s5972,s2372);
  buf x2293(s5980,s2372);
  buf x2294(s6080,s2734);
  buf x2295(s6090,s2618);
  buf x2296(s6100,s2589);
  buf x2297(s6110,s2600);
  buf x2298(s6138,s2734);
  buf x2299(s6148,s2618);
  buf x2300(s6158,s2589);
  buf x2301(s6168,s2600);
  buf x2302(s6216,s2701);
  buf x2303(s6226,s2643);
  buf x2304(s6236,s2676);
  buf x2305(s6246,s2655);
  buf x2306(s6256,s2655);
  not x2307(s6267,s6261);
  buf x2308(s6304,s2701);
  buf x2309(s6314,s2643);
  buf x2310(s6324,s2676);
  nand x2311(s6342,s6340,s6341);
  nand x2312(s6352,s6350,s6351);
  not x2313(s7351,s7345);
  not x2314(s7352,s7348);
  buf x2315(s6642,s3283);
  buf x2316(s6650,s3283);
  buf x2317(s6658,s3295);
  buf x2318(s6666,s3295);
  buf x2319(s6674,s3314);
  buf x2320(s6682,s3314);
  not x2321(s6815,s6809);
  not x2322(s6816,s6812);
  not x2323(s6825,s6819);
  not x2324(s6826,s6822);
  buf x2325(s6948,s3989);
  buf x2326(s6958,s3874);
  buf x2327(s6968,s3845);
  buf x2328(s6978,s3856);
  buf x2329(s7006,s3989);
  buf x2330(s7016,s3874);
  buf x2331(s7026,s3845);
  buf x2332(s7036,s3856);
  buf x2333(s7074,s3997);
  buf x2334(s7084,s3957);
  buf x2335(s7094,s3899);
  buf x2336(s7104,s3932);
  buf x2337(s7114,s3911);
  buf x2338(s7124,s3911);
  buf x2339(s7162,s3997);
  buf x2340(s7172,s3957);
  buf x2341(s7182,s3899);
  buf x2342(s7192,s3932);
  nand x2343(s7438,s7436,s7437);
  not x2344(s7617,s7611);
  not x2345(s7618,s7614);
  not x2346(s7609,s7603);
  not x2347(s7610,s7606);
  and x2348(s1151,s1129,s1108);
  and x2349(s1002,s902,s929);
  not x2350(s933,s929);
  and x2351(s1308,s1221,s1226,s1287);
  and x2352(s1311,s1217,s1230,s1291);
  and x2353(s1314,s1244,s1249,s1295);
  and x2354(s1317,s1240,s1253,s1299);
  and x2355(s1320,s1267,s1272,s1303);
  and x2356(s1323,s1263,s1276,s1307);
  not x2357(s1730,s1726);
  and x2358(s1789,s1702,s1726);
  and x2359(s1981,s1957,s1935);
  not x2360(s5823,s5817);
  nand x2361(s1986,s5817,s5824);
  not x2362(s5831,s5825);
  nand x2363(s1989,s5825,s5832);
  not x2364(s5839,s5833);
  nand x2365(s1993,s5833,s5840);
  not x2366(s5847,s5841);
  nand x2367(s1996,s5841,s5848);
  nand x2368(s2000,s5849,s5856);
  nand x2369(s2004,s5857,s5864);
  or x2370(s2495,s2351,s2492,s2493,s2494);
  or x2371(s2515,s2417,s2511,s2512,s2513,s2514);
  or x2372(s2757,s2597,s2754,s2755,s2756);
  or x2373(s2768,s2629,s2767);
  or x2374(s2780,s2652,s2776,s2777,s2778,s2779);
  or x2375(s2801,s2715,s2800);
  or x2376(s3046,s3028,s3045);
  or x2377(s3131,s3059,s3128,s3129,s3130);
  or x2378(s3143,s3090,s3139,s3140,s3141,s3142);
  not x2379(s3238,s3235);
  and x2380(s3258,s3216,s3235);
  or x2381(s3437,s3292,s3434,s3435,s3436);
  or x2382(s3453,s3362,s3449,s3450,s3451,s3452);
  and x2383(s3595,s3508,s3513,s3574);
  and x2384(s3598,s3504,s3517,s3578);
  or x2385(s4010,s3853,s4007,s4008,s4009);
  or x2386(s4017,s3885,s4016);
  or x2387(s4028,s3908,s4024,s4025,s4026,s4027);
  or x2388(s4048,s3971,s4047);
  and x2389(s4283,s4230,s4235,s4266);
  and x2390(s4286,s4226,s4239,s4270);
  or x2391(s4364,s4297,s4361,s4362,s4363);
  or x2392(s4376,s4324,s4372,s4373,s4374,s4375);
  and x2393(s4622,s4535,s4540,s4601);
  and x2394(s4625,s4531,s4544,s4605);
  nand x2395(s4947,s4942,s4945);
  nand x2396(s4988,s4983,s4986);
  not x2397(s5018,s5014);
  nand x2398(s5019,s5014,s5017);
  or x2399(s5024,s950,s956);
  not x2400(s5038,s5034);
  not x2401(s5106,s5102);
  nand x2402(s5107,s5102,s5105);
  not x2403(s5112,s950);
  not x2404(s5126,s5122);
  or x2405(s5468,s1715,s1749);
  not x2406(s5482,s5478);
  not x2407(s5526,s1715);
  not x2408(s5540,s5536);
  not x2409(s5588,s5584);
  nand x2410(s5589,s5584,s5587);
  or x2411(s5594,s1746,s1750);
  not x2412(s5608,s5604);
  not x2413(s5676,s5672);
  nand x2414(s5677,s5672,s5675);
  not x2415(s5682,s1746);
  not x2416(s5696,s5692);
  or x2417(s5937,s2366,s2500,s2501,s2502);
  nor x2418(s5945,s2366,s2503,s2504);
  or x2419(s5953,s2384,s2505,s2506);
  nor x2420(s5961,s2384,s2507);
  or x2421(s6070,s2612,s2762,s2763,s2764);
  nor x2422(s6128,s2612,s2765,s2766);
  nor x2423(s6264,s2693,s2798,s2799);
  nor x2424(s6284,s2670,s2792,s2793,s2794);
  nand x2425(s6360,s7348,s7351);
  nand x2426(s6361,s7345,s7352);
  or x2427(s6639,s3308,s3438,s3439,s3440);
  nor x2428(s6647,s3308,s3441,s3442);
  or x2429(s6655,s3327,s3443,s3444);
  nor x2430(s6663,s3327,s3445);
  nand x2431(s6817,s6812,s6815);
  nand x2432(s6818,s6809,s6816);
  nand x2433(s6827,s6822,s6825);
  nand x2434(s6828,s6819,s6826);
  or x2435(s6938,s3868,s4011,s4012,s4013);
  nor x2436(s6996,s3868,s4014,s4015);
  or x2437(s7044,s3949,s4042,s4043,s4044);
  or x2438(s7064,s3926,s4035,s4036,s4037,s4038);
  nor x2439(s7132,s3949,s4045,s4046);
  nor x2440(s7152,s3926,s4039,s4040,s4041);
  nand x2441(s7446,s7614,s7617);
  nand x2442(s7447,s7611,s7618);
  nand x2443(s7456,s7606,s7609);
  nand x2444(s7457,s7603,s7610);
  or x2445(s241,s1117,s1151);
  or x2446(s265,s908,s1002);
  nand x2447(s2005,s2003,s2004);
  not x2448(s4800,s4796);
  not x2449(s4808,s4804);
  not x2450(s4816,s4812);
  not x2451(s4824,s4820);
  not x2452(s4832,s4828);
  not x2453(s4848,s4844);
  not x2454(s4856,s4852);
  not x2455(s4864,s4860);
  not x2456(s4872,s4868);
  nor x2457(s1310,s1308,s1309);
  nor x2458(s1313,s1311,s1312);
  nor x2459(s1316,s1314,s1315);
  nor x2460(s1319,s1317,s1318);
  nor x2461(s1322,s1320,s1321);
  nor x2462(s1325,s1323,s1324);
  not x2463(s5392,s5388);
  or x2464(s1790,s1708,s1789);
  or x2465(s1982,s1941,s1981);
  nand x2466(s1985,s5820,s5823);
  nand x2467(s1988,s5828,s5831);
  nand x2468(s1992,s5836,s5839);
  nand x2469(s1995,s5844,s5847);
  nand x2470(s2001,s1999,s2000);
  not x2471(s2491,s2487);
  and x2472(s2508,s2420,s2472,s2436,s2409,s2454);
  and x2473(s2522,s4526,s2472,s2436,s2454,s2420);
  and x2474(s2526,s4526,s2472,s2436,s2454);
  and x2475(s2529,s4526,s2472,s2454);
  and x2476(s2531,s4526,s2472);
  not x2477(s5944,s5940);
  not x2478(s5952,s5948);
  not x2479(s5960,s5956);
  not x2480(s5968,s5964);
  nand x2481(s2555,s5972,s5975);
  not x2482(s5976,s5972);
  nand x2483(s2559,s5980,s5983);
  not x2484(s5984,s5980);
  not x2485(s2753,s2749);
  and x2486(s2771,s2742,s2701,s2676,s2655,s2643);
  and x2487(s2791,s2742,s2676,s2655,s2701);
  and x2488(s2797,s2742,s2676,s2701);
  and x2489(s2807,s2742,s2701);
  not x2490(s6114,s6110);
  not x2491(s6172,s6168);
  not x2492(s6250,s6246);
  not x2493(s6260,s6256);
  not x2494(s6346,s6342);
  not x2495(s6356,s6352);
  not x2496(s3127,s3123);
  and x2497(s3156,s3123,s3136);
  or x2498(s3259,s3223,s3258);
  and x2499(s3466,s3431,s3446);
  not x2500(s6646,s6642);
  not x2501(s6654,s6650);
  not x2502(s6662,s6658);
  not x2503(s6670,s6666);
  nand x2504(s3483,s6674,s6677);
  not x2505(s6678,s6674);
  nand x2506(s3487,s6682,s6685);
  not x2507(s6686,s6682);
  not x2508(s3582,s3579);
  not x2509(s3586,s3583);
  not x2510(s3590,s3587);
  not x2511(s3594,s3591);
  nor x2512(s3597,s3595,s3596);
  nor x2513(s3600,s3598,s3599);
  and x2514(s3602,s3536,s3527,s3579);
  and x2515(s3605,s3540,s3531,s3583);
  and x2516(s3608,s3559,s3550,s3587);
  and x2517(s3611,s3563,s3554,s3591);
  not x2518(s4023,s4020);
  not x2519(s6982,s6978);
  not x2520(s7040,s7036);
  not x2521(s7118,s7114);
  not x2522(s7128,s7124);
  and x2523(s4089,s4004,s4020);
  not x2524(s4250,s4247);
  not x2525(s4254,s4251);
  not x2526(s4258,s4255);
  not x2527(s4262,s4259);
  and x2528(s4272,s4189,s4180,s4247);
  and x2529(s4275,s4193,s4184,s4251);
  and x2530(s4278,s4212,s4203,s4255);
  and x2531(s4281,s4216,s4207,s4259);
  nor x2532(s4285,s4283,s4284);
  nor x2533(s4288,s4286,s4287);
  not x2534(s4360,s4356);
  nand x2535(s4380,s4369,s89);
  and x2536(s4386,s4356,s4369);
  not x2537(s7442,s7438);
  not x2538(s4609,s4606);
  not x2539(s4613,s4610);
  not x2540(s4617,s4614);
  not x2541(s4621,s4618);
  nor x2542(s4624,s4622,s4623);
  nor x2543(s4627,s4625,s4626);
  and x2544(s4629,s4563,s4554,s4606);
  and x2545(s4632,s4567,s4558,s4610);
  and x2546(s4635,s4586,s4577,s4614);
  and x2547(s4638,s4590,s4581,s4618);
  buf x2548(s4836,s2472);
  nand x2549(s4949,s4947,s4948);
  nand x2550(s4990,s4988,s4989);
  nand x2551(s5020,s5011,s5018);
  nand x2552(s5108,s5099,s5106);
  nand x2553(s5590,s5581,s5588);
  nand x2554(s5678,s5669,s5676);
  not x2555(s6084,s6080);
  not x2556(s6094,s6090);
  not x2557(s6104,s6100);
  not x2558(s6142,s6138);
  not x2559(s6152,s6148);
  not x2560(s6162,s6158);
  buf x2561(s6206,s2742);
  not x2562(s6220,s6216);
  not x2563(s6230,s6226);
  not x2564(s6240,s6236);
  not x2565(s6328,s6324);
  buf x2566(s6294,s2742);
  not x2567(s6308,s6304);
  not x2568(s6318,s6314);
  nand x2569(s6362,s6360,s6361);
  nand x2570(s6840,s6817,s6818);
  nand x2571(s6848,s6827,s6828);
  not x2572(s6952,s6948);
  not x2573(s6962,s6958);
  not x2574(s6972,s6968);
  not x2575(s7010,s7006);
  not x2576(s7020,s7016);
  not x2577(s7030,s7026);
  not x2578(s7078,s7074);
  not x2579(s7088,s7084);
  not x2580(s7098,s7094);
  not x2581(s7108,s7104);
  not x2582(s7196,s7192);
  not x2583(s7166,s7162);
  not x2584(s7176,s7172);
  not x2585(s7186,s7182);
  nand x2586(s7448,s7446,s7447);
  nand x2587(s7458,s7456,s7457);
  and x2588(s254,s3046,s3249);
  and x2589(s260,s3046,s3249);
  nand x2590(s1987,s1985,s1986);
  nand x2591(s1994,s1992,s1993);
  not x2592(s2002,s2001);
  and x2593(s962,s933,s924);
  and x2594(s1751,s1730,s1721);
  nand x2595(s1990,s1988,s1989);
  nand x2596(s1997,s1995,s1996);
  not x2597(s2499,s2495);
  and x2598(s2536,s2515,s2487);
  not x2599(s5943,s5937);
  nand x2600(s2542,s5937,s5944);
  not x2601(s5951,s5945);
  nand x2602(s2545,s5945,s5952);
  not x2603(s5959,s5953);
  nand x2604(s2549,s5953,s5960);
  not x2605(s5967,s5961);
  nand x2606(s2552,s5961,s5968);
  nand x2607(s2556,s5969,s5976);
  nand x2608(s2560,s5977,s5984);
  not x2609(s2761,s2757);
  not x2610(s2784,s2780);
  and x2611(s2853,s2749,s2780);
  not x2612(s3135,s3131);
  not x2613(s3146,s3143);
  and x2614(s3163,s3123,s3143);
  and x2615(s3467,s3453,s3431);
  not x2616(s6645,s6639);
  nand x2617(s3470,s6639,s6646);
  not x2618(s6653,s6647);
  nand x2619(s3473,s6647,s6654);
  not x2620(s6661,s6655);
  nand x2621(s3477,s6655,s6662);
  not x2622(s6669,s6663);
  nand x2623(s3480,s6663,s6670);
  nand x2624(s3484,s6671,s6678);
  nand x2625(s3488,s6679,s6686);
  and x2626(s3601,s3531,s3536,s3582);
  and x2627(s3604,s3527,s3540,s3586);
  and x2628(s3607,s3554,s3559,s3590);
  and x2629(s3610,s3550,s3563,s3594);
  not x2630(s4032,s4028);
  and x2631(s4090,s4004,s4028);
  and x2632(s4271,s4184,s4189,s4250);
  and x2633(s4274,s4180,s4193,s4254);
  and x2634(s4277,s4207,s4212,s4258);
  and x2635(s4280,s4203,s4216,s4262);
  not x2636(s4368,s4364);
  not x2637(s4379,s4376);
  and x2638(s4387,s4356,s4376);
  and x2639(s4628,s4558,s4563,s4609);
  and x2640(s4631,s4554,s4567,s4613);
  and x2641(s4634,s4581,s4586,s4617);
  and x2642(s4637,s4577,s4590,s4621);
  or x2643(s4841,s2431,s2518,s2519,s2520,s2522);
  or x2644(s4849,s2448,s2523,s2524,s2526);
  or x2645(s4857,s2465,s2527,s2529);
  or x2646(s4865,s2481,s2531);
  nand x2647(s5021,s5019,s5020);
  not x2648(s5028,s5024);
  nand x2649(s5109,s5107,s5108);
  not x2650(s5116,s5112);
  nand x2651(s5369,s1313,s1310);
  nand x2652(s5377,s1319,s1316);
  nand x2653(s5385,s1325,s1322);
  not x2654(s5472,s5468);
  nand x2655(s5473,s5468,s5471);
  not x2656(s5530,s5526);
  nand x2657(s5531,s5526,s5529);
  nand x2658(s5591,s5589,s5590);
  not x2659(s5598,s5594);
  nand x2660(s5679,s5677,s5678);
  not x2661(s5686,s5682);
  or x2662(s6060,s2768,s2804);
  not x2663(s6074,s6070);
  not x2664(s6118,s2768);
  not x2665(s6132,s6128);
  or x2666(s6176,s2693,s2795,s2796,s2797);
  or x2667(s6186,s2801,s2807);
  or x2668(s6196,s2670,s2788,s2789,s2790,s2791);
  not x2669(s6268,s6264);
  nand x2670(s6269,s6264,s6267);
  not x2671(s6274,s2801);
  not x2672(s6288,s6284);
  nand x2673(s6337,s4288,s4285);
  nand x2674(s6829,s3600,s3597);
  or x2675(s6928,s4017,s4051);
  not x2676(s6942,s6938);
  not x2677(s6986,s4017);
  not x2678(s7000,s6996);
  not x2679(s7048,s7044);
  nand x2680(s7049,s7044,s7047);
  or x2681(s7054,s4048,s4052);
  not x2682(s7068,s7064);
  not x2683(s7136,s7132);
  nand x2684(s7137,s7132,s7135);
  not x2685(s7142,s4048);
  not x2686(s7156,s7152);
  nand x2687(s7433,s4627,s4624);
  and x2688(s242,s1982,s1146);
  nand x2689(s3151,s3135,s3127);
  and x2690(s257,s89,s4386,s3156,s3035,s3249);
  and x2691(s263,s89,s4386,s3156,s3035,s3249);
  and x2692(s266,s1790,s997);
  not x2693(s1991,s1990);
  not x2694(s1998,s1997);
  nand x2695(s3489,s3487,s3488);
  nand x2696(s371,s4836,s4839);
  not x2697(s4840,s4836);
  nand x2698(s2561,s2559,s2560);
  and x2699(s2532,s2487,s2508);
  or x2700(s2537,s2495,s2536);
  nand x2701(s2541,s5940,s5943);
  nand x2702(s2544,s5948,s5951);
  nand x2703(s2548,s5956,s5959);
  nand x2704(s2551,s5964,s5967);
  nand x2705(s2557,s2555,s2556);
  and x2706(s2563,s2508,s4526);
  nand x2707(s2577,s2499,s2491);
  not x2708(s2775,s2771);
  nand x2709(s2806,s2771,s4526);
  nand x2710(s2808,s2761,s2753);
  and x2711(s2852,s2749,s2771);
  or x2712(s2854,s2757,s2853);
  not x2713(s6366,s6362);
  nand x2714(s4381,s4368,s4360);
  or x2715(s3164,s3131,s3163);
  and x2716(s3241,s89,s4386,s3156,s3035);
  or x2717(s3468,s3437,s3467);
  nand x2718(s3469,s6642,s6645);
  nand x2719(s3472,s6650,s6653);
  nand x2720(s3476,s6658,s6661);
  nand x2721(s3479,s6666,s6669);
  nand x2722(s3485,s3483,s3484);
  nor x2723(s3603,s3601,s3602);
  nor x2724(s3606,s3604,s3605);
  nor x2725(s3609,s3607,s3608);
  nor x2726(s3612,s3610,s3611);
  not x2727(s6844,s6840);
  not x2728(s6852,s6848);
  or x2729(s4091,s4010,s4090);
  nor x2730(s4273,s4271,s4272);
  nor x2731(s4276,s4274,s4275);
  nor x2732(s4279,s4277,s4278);
  nor x2733(s4282,s4280,s4281);
  and x2734(s4382,s4379,s4380);
  or x2735(s4388,s4364,s4387);
  not x2736(s7452,s7448);
  not x2737(s7462,s7458);
  nor x2738(s4630,s4628,s4629);
  nor x2739(s4633,s4631,s4632);
  nor x2740(s4636,s4634,s4635);
  nor x2741(s4639,s4637,s4638);
  not x2742(s4955,s4949);
  nand x2743(s4958,s4949,s4956);
  not x2744(s4996,s4990);
  nand x2745(s4999,s4990,s4997);
  nand x2746(s5474,s5465,s5472);
  nand x2747(s5532,s5523,s5530);
  not x2748(s6210,s6206);
  nand x2749(s6270,s6261,s6268);
  not x2750(s6298,s6294);
  nand x2751(s7050,s7041,s7048);
  nand x2752(s7138,s7129,s7136);
  nand x2753(s3471,s3469,s3470);
  nand x2754(s3478,s3476,s3477);
  not x2755(s3486,s3485);
  nand x2756(s372,s4833,s4840);
  nand x2757(s2543,s2541,s2542);
  nand x2758(s2550,s2548,s2549);
  not x2759(s2558,s2557);
  not x2760(s4847,s4841);
  nand x2761(s387,s4841,s4848);
  not x2762(s4855,s4849);
  nand x2763(s390,s4849,s4856);
  not x2764(s4863,s4857);
  nand x2765(s393,s4857,s4864);
  not x2766(s4871,s4865);
  nand x2767(s396,s4865,s4872);
  not x2768(s965,s962);
  not x2769(s5375,s5369);
  nand x2770(s1327,s5369,s5376);
  not x2771(s5383,s5377);
  nand x2772(s1330,s5377,s5384);
  not x2773(s5391,s5385);
  nand x2774(s1333,s5385,s5392);
  not x2775(s1754,s1751);
  nand x2776(s2546,s2544,s2545);
  nand x2777(s2553,s2551,s2552);
  or x2778(s2564,s2515,s2563);
  and x2779(s2809,s2784,s2806);
  and x2780(s2813,s2784,s2775);
  not x2781(s6345,s6337);
  nand x2782(s2860,s6337,s6346);
  nand x2783(s3474,s3472,s3473);
  nand x2784(s3481,s3479,s3480);
  not x2785(s6835,s6829);
  nand x2786(s3614,s6829,s6836);
  and x2787(s4053,s4032,s4023);
  not x2788(s7441,s7433);
  nand x2789(s4516,s7433,s7442);
  nand x2790(s4957,s4952,s4955);
  nand x2791(s4998,s4993,s4996);
  not x2792(s5027,s5021);
  nand x2793(s5030,s5021,s5028);
  not x2794(s5115,s5109);
  nand x2795(s5118,s5109,s5116);
  nand x2796(s5475,s5473,s5474);
  nand x2797(s5533,s5531,s5532);
  not x2798(s5597,s5591);
  nand x2799(s5600,s5591,s5598);
  not x2800(s5685,s5679);
  nand x2801(s5688,s5679,s5686);
  not x2802(s6064,s6060);
  nand x2803(s6065,s6060,s6063);
  not x2804(s6122,s6118);
  nand x2805(s6123,s6118,s6121);
  not x2806(s6180,s6176);
  nand x2807(s6181,s6176,s6179);
  not x2808(s6190,s6186);
  not x2809(s6200,s6196);
  nand x2810(s6271,s6269,s6270);
  not x2811(s6278,s6274);
  nand x2812(s6347,s4276,s4273);
  nand x2813(s6357,s4282,s4279);
  nand x2814(s6837,s3606,s3603);
  nand x2815(s6845,s3612,s3609);
  not x2816(s6932,s6928);
  nand x2817(s6933,s6928,s6931);
  not x2818(s6990,s6986);
  nand x2819(s6991,s6986,s6989);
  nand x2820(s7051,s7049,s7050);
  not x2821(s7058,s7054);
  nand x2822(s7139,s7137,s7138);
  not x2823(s7146,s7142);
  nand x2824(s7443,s4639,s4636);
  nand x2825(s7453,s4633,s4630);
  and x2826(s243,s3468,s1974,s1146);
  and x2827(s244,s2537,s3466,s1974,s1146);
  and x2828(s245,s4526,s2532,s3466,s1974,s1146);
  and x2829(s255,s3164,s3035,s3249);
  and x2830(s256,s4388,s3156,s3035,s3249);
  and x2831(s261,s3164,s3035,s3249);
  and x2832(s262,s4388,s3156,s3035,s3249);
  and x2833(s267,s4091,s1788,s997);
  and x2834(s268,s2854,s4089,s1788,s997);
  and x2835(s269,s4526,s2852,s4089,s1788,s997);
  not x2836(s3475,s3474);
  not x2837(s3482,s3481);
  nand x2838(s373,s371,s372);
  not x2839(s2547,s2546);
  not x2840(s2554,s2553);
  nand x2841(s386,s4844,s4847);
  nand x2842(s389,s4852,s4855);
  nand x2843(s392,s4860,s4863);
  nand x2844(s395,s4868,s4871);
  nand x2845(s1326,s5372,s5375);
  nand x2846(s1329,s5380,s5383);
  nand x2847(s1332,s5388,s5391);
  and x2848(s1436,s4091,s1788);
  and x2849(s1440,s2854,s4089,s1788);
  and x2850(s1445,s4526,s2852,s4089,s1788);
  and x2851(s1450,s2854,s4089);
  and x2852(s1454,s4526,s2852,s4089);
  nand x2853(s2859,s6342,s6345);
  not x2854(s4385,s4382);
  and x2855(s3148,s4382,s4364);
  and x2856(s3239,s3164,s3035);
  and x2857(s3240,s4388,s3156,s3035);
  and x2858(s3265,s3468,s1974);
  and x2859(s3267,s2537,s3466,s1974);
  and x2860(s3270,s4526,s2532,s3466,s1974);
  and x2861(s3274,s2537,s3466);
  and x2862(s3277,s4526,s2532,s3466);
  nand x2863(s3613,s6832,s6835);
  nand x2864(s4515,s7438,s7441);
  nand x2865(s4959,s4957,s4958);
  nand x2866(s5000,s4998,s4999);
  nand x2867(s5029,s5024,s5027);
  nand x2868(s5117,s5112,s5115);
  nand x2869(s5599,s5594,s5597);
  nand x2870(s5687,s5682,s5685);
  nand x2871(s6066,s6057,s6064);
  nand x2872(s6124,s6115,s6122);
  nand x2873(s6182,s6173,s6180);
  nand x2874(s6934,s6925,s6932);
  nand x2875(s6992,s6983,s6990);
  or x2876(s246,s241,s242,s243,s244,s245);
  or x2877(s258,s3259,s254,s255,s256,s257);
  or x2878(s264,s3259,s260,s261,s262,s263);
  or x2879(s270,s265,s266,s267,s268,s269);
  and x2880(s375,s2564,s2543);
  and x2881(s378,s2564,s2550);
  and x2882(s381,s2564,s2558);
  and x2883(s384,s2564,s2406);
  nand x2884(s388,s386,s387);
  nand x2885(s391,s389,s390);
  nand x2886(s394,s392,s393);
  nand x2887(s397,s395,s396);
  nand x2888(s1328,s1326,s1327);
  nand x2889(s1331,s1329,s1330);
  nand x2890(s1334,s1332,s1333);
  or x2891(s1447,s1790,s1436,s1440,s1445);
  or x2892(s1766,s4091,s1450,s1454);
  not x2893(s2571,s2564);
  and x2894(s2579,s2577,s2564);
  not x2895(s2812,s2809);
  not x2896(s2816,s2813);
  and x2897(s2851,s2809,s2757);
  nand x2898(s2861,s2859,s2860);
  not x2899(s6355,s6347);
  nand x2900(s2863,s6347,s6356);
  not x2901(s6365,s6357);
  nand x2902(s2866,s6357,s6366);
  and x2903(s3147,s4381,s4385);
  or x2904(s3242,s3046,s3239,s3240,s3241);
  or x2905(s3271,s1982,s3265,s3267,s3270);
  or x2906(s3279,s3468,s3274,s3277);
  nand x2907(s3615,s3613,s3614);
  not x2908(s6843,s6837);
  nand x2909(s3617,s6837,s6844);
  not x2910(s6851,s6845);
  nand x2911(s3620,s6845,s6852);
  not x2912(s4056,s4053);
  nand x2913(s4517,s4515,s4516);
  not x2914(s7451,s7443);
  nand x2915(s4519,s7443,s7452);
  not x2916(s7461,s7453);
  nand x2917(s4522,s7453,s7462);
  nand x2918(s5031,s5029,s5030);
  nand x2919(s5119,s5117,s5118);
  not x2920(s5481,s5475);
  nand x2921(s5484,s5475,s5482);
  not x2922(s5539,s5533);
  nand x2923(s5542,s5533,s5540);
  nand x2924(s5601,s5599,s5600);
  nand x2925(s5689,s5687,s5688);
  nand x2926(s6067,s6065,s6066);
  nand x2927(s6125,s6123,s6124);
  nand x2928(s6183,s6181,s6182);
  not x2929(s6277,s6271);
  nand x2930(s6280,s6271,s6278);
  nand x2931(s6935,s6933,s6934);
  nand x2932(s6993,s6991,s6992);
  not x2933(s7057,s7051);
  nand x2934(s7060,s7051,s7058);
  not x2935(s7145,s7139);
  nand x2936(s7148,s7139,s7146);
  nand x2937(s4968,s4959,s4966);
  nand x2938(s5009,s5000,s5007);
  and x2939(s2850,s2808,s2812);
  nand x2940(s2862,s6352,s6355);
  nand x2941(s2865,s6362,s6365);
  or x2942(s3149,s3147,s3148);
  nand x2943(s3243,s3228,s3242);
  nand x2944(s3616,s6840,s6843);
  nand x2945(s3619,s6848,s6851);
  nand x2946(s4518,s7448,s7451);
  nand x2947(s4521,s7458,s7461);
  not x2948(s4965,s4959);
  not x2949(s5006,s5000);
  nand x2950(s5483,s5478,s5481);
  nand x2951(s5541,s5536,s5539);
  nand x2952(s6279,s6274,s6277);
  nand x2953(s7059,s7054,s7057);
  nand x2954(s7147,s7142,s7145);
  and x2955(s374,s2547,s2571);
  and x2956(s377,s2554,s2571);
  and x2957(s380,s2561,s2571);
  and x2958(s383,s2400,s2571);
  nand x2959(s955,s920,s1447);
  nand x2960(s4967,s4962,s4965);
  nand x2961(s5008,s5003,s5006);
  buf x2962(s975,s1447);
  and x2963(s1136,s3271,s1093,s1055,s1074,s1038);
  and x2964(s1140,s3271,s1093,s1055,s1074);
  and x2965(s1143,s3271,s1093,s1074);
  and x2966(s1145,s3271,s1093);
  and x2967(s1160,s1122,s3271);
  not x2968(s1771,s1766);
  and x2969(s1964,s3279,s1921,s1885,s1903,s1869);
  and x2970(s1968,s3279,s1921,s1885,s1903);
  and x2971(s1971,s3279,s1921,s1903);
  and x2972(s1973,s3279,s1921);
  and x2973(s2007,s1950,s3279);
  and x2974(s2578,s2495,s2571);
  nand x2975(s2864,s2862,s2863);
  nand x2976(s2867,s2865,s2866);
  nand x2977(s3150,s3136,s3149);
  and x2978(s3245,s3238,s3243);
  nand x2979(s3618,s3616,s3617);
  nand x2980(s3621,s3619,s3620);
  or x2981(s4067,s2850,s2851);
  nand x2982(s4520,s4518,s4519);
  nand x2983(s4523,s4521,s4522);
  buf x2984(s4713,s3279);
  buf x2985(s4753,s3271);
  not x2986(s5037,s5031);
  nand x2987(s5040,s5031,s5038);
  not x2988(s5125,s5119);
  nand x2989(s5128,s5119,s5126);
  nand x2990(s5485,s5483,s5484);
  nand x2991(s5543,s5541,s5542);
  not x2992(s5607,s5601);
  nand x2993(s5610,s5601,s5608);
  not x2994(s5695,s5689);
  nand x2995(s5698,s5689,s5696);
  not x2996(s6073,s6067);
  nand x2997(s6076,s6067,s6074);
  not x2998(s6131,s6125);
  nand x2999(s6134,s6125,s6132);
  not x3000(s6189,s6183);
  nand x3001(s6192,s6183,s6190);
  nand x3002(s6281,s6279,s6280);
  not x3003(s6941,s6935);
  nand x3004(s6944,s6935,s6942);
  not x3005(s6999,s6993);
  nand x3006(s7002,s6993,s7000);
  nand x3007(s7061,s7059,s7060);
  nand x3008(s7149,s7147,s7148);
  or x3009(s376,s374,s375);
  or x3010(s379,s377,s378);
  or x3011(s382,s380,s381);
  or x3012(s385,s383,s384);
  and x3013(s958,s933,s955);
  nand x3014(s967,s4967,s4968);
  nand x3015(s971,s5008,s5009);
  or x3016(s1161,s1129,s1160);
  or x3017(s2008,s1957,s2007);
  or x3018(s2580,s2578,s2579);
  and x3019(s2868,s1331,s2861,s2864,s2867);
  and x3020(s3152,s3146,s3150);
  and x3021(s4443,s1328,s1334,s3618,s3621);
  and x3022(s4524,s3615,s4517,s4520,s4523);
  or x3023(s4721,s1880,s1960,s1961,s1962,s1964);
  or x3024(s4729,s1897,s1965,s1966,s1968);
  or x3025(s4737,s1914,s1969,s1971);
  or x3026(s4745,s1929,s1973);
  or x3027(s4761,s1050,s1132,s1133,s1134,s1136);
  or x3028(s4769,s1068,s1137,s1138,s1140);
  or x3029(s4777,s1086,s1141,s1143);
  or x3030(s4785,s1102,s1145);
  nand x3031(s5039,s5034,s5037);
  nand x3032(s5127,s5122,s5125);
  nand x3033(s5609,s5604,s5607);
  nand x3034(s5697,s5692,s5695);
  nand x3035(s6075,s6070,s6073);
  nand x3036(s6133,s6128,s6131);
  nand x3037(s6191,s6186,s6189);
  nand x3038(s6943,s6938,s6941);
  nand x3039(s7001,s6996,s6999);
  not x3040(s3248,s3245);
  and x3041(s248,s3245,s3223);
  not x3042(s4719,s4713);
  nand x3043(s294,s4713,s4720);
  not x3044(s4759,s4753);
  nand x3045(s323,s4753,s4760);
  not x3046(s980,s975);
  not x3047(s4072,s4067);
  nand x3048(s5041,s5039,s5040);
  nand x3049(s5129,s5127,s5128);
  not x3050(s5491,s5485);
  nand x3051(s5494,s5485,s5492);
  not x3052(s5549,s5543);
  nand x3053(s5552,s5543,s5550);
  nand x3054(s5611,s5609,s5610);
  nand x3055(s5699,s5697,s5698);
  nand x3056(s6077,s6075,s6076);
  nand x3057(s6135,s6133,s6134);
  nand x3058(s6193,s6191,s6192);
  not x3059(s6287,s6281);
  nand x3060(s6290,s6281,s6288);
  nand x3061(s6945,s6943,s6944);
  nand x3062(s7003,s7001,s7002);
  not x3063(s7067,s7061);
  nand x3064(s7070,s7061,s7068);
  not x3065(s7155,s7149);
  nand x3066(s7158,s7149,s7156);
  and x3067(s247,s3244,s3248);
  not x3068(s3155,s3152);
  and x3069(s251,s3152,s3131);
  and x3070(s272,s1176,s1161);
  not x3071(s961,s958);
  and x3072(s275,s958,s908);
  nand x3073(s293,s4716,s4719);
  and x3074(s297,s2008,s1987);
  and x3075(s300,s2008,s1994);
  and x3076(s303,s2008,s2002);
  and x3077(s306,s2008,s1856);
  not x3078(s4727,s4721);
  nand x3079(s309,s4721,s4728);
  not x3080(s4735,s4729);
  nand x3081(s312,s4729,s4736);
  not x3082(s4743,s4737);
  nand x3083(s315,s4737,s4744);
  not x3084(s4751,s4745);
  nand x3085(s318,s4745,s4752);
  nand x3086(s322,s4756,s4759);
  not x3087(s4767,s4761);
  nand x3088(s326,s4761,s4768);
  not x3089(s4775,s4769);
  nand x3090(s329,s4769,s4776);
  not x3091(s4783,s4777);
  nand x3092(s332,s4777,s4784);
  not x3093(s4791,s4785);
  nand x3094(s335,s4785,s4792);
  not x3095(s412,s4443);
  not x3096(s414,s4524);
  not x3097(s416,s2868);
  and x3098(s2881,s4443,s4524,s2868);
  and x3099(s993,s971,s962,s975);
  and x3100(s994,s967,s965,s975);
  not x3101(s1166,s1161);
  and x3102(s1171,s1161,s1155);
  and x3103(s1174,s1161,s1023);
  not x3104(s2014,s2008);
  and x3105(s3459,s2580,s3417,s3381,s3399,s3365);
  and x3106(s3462,s2580,s3417,s3381,s3399);
  and x3107(s3464,s2580,s3417,s3399);
  and x3108(s3465,s2580,s3417);
  and x3109(s3490,s3446,s2580);
  buf x3110(s4793,s2580);
  nand x3111(s5493,s5488,s5491);
  nand x3112(s5551,s5546,s5549);
  nand x3113(s6289,s6284,s6287);
  nand x3114(s7069,s7064,s7067);
  nand x3115(s7157,s7152,s7155);
  or x3116(s249,s247,s248);
  and x3117(s250,s3151,s3155);
  and x3118(s274,s957,s961);
  nand x3119(s295,s293,s294);
  nand x3120(s308,s4724,s4727);
  nand x3121(s311,s4732,s4735);
  nand x3122(s314,s4740,s4743);
  nand x3123(s317,s4748,s4751);
  nand x3124(s324,s322,s323);
  nand x3125(s325,s4764,s4767);
  nand x3126(s328,s4772,s4775);
  nand x3127(s331,s4780,s4783);
  nand x3128(s334,s4788,s4791);
  and x3129(s417,s2876,s2878,s2881);
  and x3130(s991,s971,s933,s980);
  and x3131(s992,s967,s929,s980);
  or x3132(s3491,s3453,s3490);
  or x3133(s4801,s3376,s3456,s3457,s3458,s3459);
  or x3134(s4809,s3393,s3460,s3461,s3462);
  or x3135(s4817,s3410,s3463,s3464);
  or x3136(s4825,s3425,s3465);
  not x3137(s5047,s5041);
  nand x3138(s5050,s5041,s5048);
  not x3139(s5135,s5129);
  nand x3140(s5138,s5129,s5136);
  nand x3141(s5495,s5493,s5494);
  nand x3142(s5553,s5551,s5552);
  not x3143(s5617,s5611);
  nand x3144(s5620,s5611,s5618);
  not x3145(s5705,s5699);
  nand x3146(s5708,s5699,s5706);
  not x3147(s6083,s6077);
  nand x3148(s6086,s6077,s6084);
  not x3149(s6141,s6135);
  nand x3150(s6144,s6135,s6142);
  not x3151(s6199,s6193);
  nand x3152(s6202,s6193,s6200);
  nand x3153(s6291,s6289,s6290);
  not x3154(s6951,s6945);
  nand x3155(s6954,s6945,s6952);
  not x3156(s7009,s7003);
  nand x3157(s7012,s7003,s7010);
  nand x3158(s7071,s7069,s7070);
  nand x3159(s7159,s7157,s7158);
  or x3160(s252,s250,s251);
  and x3161(s271,s1117,s1166);
  or x3162(s276,s274,s275);
  and x3163(s296,s1991,s2014);
  and x3164(s299,s1998,s2014);
  and x3165(s302,s2005,s2014);
  and x3166(s305,s1850,s2014);
  nand x3167(s310,s308,s309);
  nand x3168(s313,s311,s312);
  nand x3169(s316,s314,s315);
  nand x3170(s319,s317,s318);
  nand x3171(s327,s325,s326);
  nand x3172(s330,s328,s329);
  nand x3173(s333,s331,s332);
  nand x3174(s336,s334,s335);
  not x3175(s4799,s4793);
  nand x3176(s343,s4793,s4800);
  not x3177(s418,s417);
  and x3178(s1170,s1158,s1166);
  and x3179(s1173,s1019,s1166);
  nand x3180(s5049,s5044,s5047);
  nand x3181(s5137,s5132,s5135);
  or x3182(s5167,s991,s992,s993,s994);
  nand x3183(s5619,s5614,s5617);
  nand x3184(s5707,s5702,s5705);
  nand x3185(s6085,s6080,s6083);
  nand x3186(s6143,s6138,s6141);
  nand x3187(s6201,s6196,s6199);
  nand x3188(s6953,s6948,s6951);
  nand x3189(s7011,s7006,s7009);
  or x3190(s273,s271,s272);
  or x3191(s298,s296,s297);
  or x3192(s301,s299,s300);
  or x3193(s304,s302,s303);
  or x3194(s307,s305,s306);
  nand x3195(s342,s4796,s4799);
  and x3196(s346,s3491,s3471);
  and x3197(s349,s3491,s3478);
  and x3198(s352,s3491,s3486);
  and x3199(s355,s3491,s3350);
  not x3200(s4807,s4801);
  nand x3201(s358,s4801,s4808);
  not x3202(s4815,s4809);
  nand x3203(s361,s4809,s4816);
  not x3204(s4823,s4817);
  nand x3205(s364,s4817,s4824);
  not x3206(s4831,s4825);
  nand x3207(s367,s4825,s4832);
  or x3208(s1172,s1170,s1171);
  or x3209(s1175,s1173,s1174);
  not x3210(s3497,s3491);
  nand x3211(s5051,s5049,s5050);
  nand x3212(s5139,s5137,s5138);
  not x3213(s5501,s5495);
  nand x3214(s5504,s5495,s5502);
  not x3215(s5559,s5553);
  nand x3216(s5562,s5553,s5560);
  nand x3217(s5621,s5619,s5620);
  nand x3218(s5709,s5707,s5708);
  nand x3219(s6087,s6085,s6086);
  nand x3220(s6145,s6143,s6144);
  nand x3221(s6203,s6201,s6202);
  not x3222(s6297,s6291);
  nand x3223(s6300,s6291,s6298);
  nand x3224(s6955,s6953,s6954);
  nand x3225(s7013,s7011,s7012);
  not x3226(s7077,s7071);
  nand x3227(s7080,s7071,s7078);
  not x3228(s7165,s7159);
  nand x3229(s7168,s7159,s7166);
  nand x3230(s344,s342,s343);
  nand x3231(s357,s4804,s4807);
  nand x3232(s360,s4812,s4815);
  nand x3233(s363,s4820,s4823);
  nand x3234(s366,s4828,s4831);
  not x3235(s5173,s5167);
  buf x3236(s422,s1172);
  buf x3237(s469,s1172);
  buf x3238(s419,s1175);
  buf x3239(s471,s1175);
  nand x3240(s5503,s5498,s5501);
  nand x3241(s5561,s5556,s5559);
  nand x3242(s6299,s6294,s6297);
  nand x3243(s7079,s7074,s7077);
  nand x3244(s7167,s7162,s7165);
  and x3245(s345,s3475,s3497);
  and x3246(s348,s3482,s3497);
  and x3247(s351,s3489,s3497);
  and x3248(s354,s3344,s3497);
  nand x3249(s359,s357,s358);
  nand x3250(s362,s360,s361);
  nand x3251(s365,s363,s364);
  nand x3252(s368,s366,s367);
  not x3253(s5057,s5051);
  nand x3254(s5060,s5051,s5058);
  not x3255(s5145,s5139);
  nand x3256(s5148,s5139,s5146);
  nand x3257(s5505,s5503,s5504);
  nand x3258(s5563,s5561,s5562);
  not x3259(s5627,s5621);
  nand x3260(s5630,s5621,s5628);
  not x3261(s5715,s5709);
  nand x3262(s5718,s5709,s5716);
  not x3263(s6093,s6087);
  nand x3264(s6096,s6087,s6094);
  not x3265(s6151,s6145);
  nand x3266(s6154,s6145,s6152);
  not x3267(s6209,s6203);
  nand x3268(s6212,s6203,s6210);
  nand x3269(s6301,s6299,s6300);
  not x3270(s6961,s6955);
  nand x3271(s6964,s6955,s6962);
  not x3272(s7019,s7013);
  nand x3273(s7022,s7013,s7020);
  nand x3274(s7081,s7079,s7080);
  nand x3275(s7169,s7167,s7168);
  or x3276(s347,s345,s346);
  or x3277(s350,s348,s349);
  or x3278(s353,s351,s352);
  or x3279(s356,s354,s355);
  nand x3280(s5059,s5054,s5057);
  nand x3281(s5147,s5142,s5145);
  nand x3282(s5629,s5624,s5627);
  nand x3283(s5717,s5712,s5715);
  nand x3284(s6095,s6090,s6093);
  nand x3285(s6153,s6148,s6151);
  nand x3286(s6211,s6206,s6209);
  nand x3287(s6963,s6958,s6961);
  nand x3288(s7021,s7016,s7019);
  nand x3289(s5061,s5059,s5060);
  nand x3290(s5149,s5147,s5148);
  not x3291(s5511,s5505);
  nand x3292(s5514,s5505,s5512);
  not x3293(s5569,s5563);
  nand x3294(s5572,s5563,s5570);
  nand x3295(s5631,s5629,s5630);
  nand x3296(s5719,s5717,s5718);
  nand x3297(s6097,s6095,s6096);
  nand x3298(s6155,s6153,s6154);
  nand x3299(s6213,s6211,s6212);
  not x3300(s6307,s6301);
  nand x3301(s6310,s6301,s6308);
  nand x3302(s6965,s6963,s6964);
  nand x3303(s7023,s7021,s7022);
  not x3304(s7087,s7081);
  nand x3305(s7090,s7081,s7088);
  not x3306(s7175,s7169);
  nand x3307(s7178,s7169,s7176);
  nand x3308(s5513,s5508,s5511);
  nand x3309(s5571,s5566,s5569);
  nand x3310(s6309,s6304,s6307);
  nand x3311(s7089,s7084,s7087);
  nand x3312(s7177,s7172,s7175);
  not x3313(s5067,s5061);
  nand x3314(s5070,s5061,s5068);
  not x3315(s5155,s5149);
  nand x3316(s5158,s5149,s5156);
  nand x3317(s5515,s5513,s5514);
  nand x3318(s5573,s5571,s5572);
  not x3319(s5637,s5631);
  nand x3320(s5640,s5631,s5638);
  not x3321(s5725,s5719);
  nand x3322(s5728,s5719,s5726);
  not x3323(s6103,s6097);
  nand x3324(s6106,s6097,s6104);
  not x3325(s6161,s6155);
  nand x3326(s6164,s6155,s6162);
  not x3327(s6219,s6213);
  nand x3328(s6222,s6213,s6220);
  nand x3329(s6311,s6309,s6310);
  not x3330(s6971,s6965);
  nand x3331(s6974,s6965,s6972);
  not x3332(s7029,s7023);
  nand x3333(s7032,s7023,s7030);
  nand x3334(s7091,s7089,s7090);
  nand x3335(s7179,s7177,s7178);
  nand x3336(s5069,s5064,s5067);
  nand x3337(s5157,s5152,s5155);
  nand x3338(s5639,s5634,s5637);
  nand x3339(s5727,s5722,s5725);
  nand x3340(s6105,s6100,s6103);
  nand x3341(s6163,s6158,s6161);
  nand x3342(s6221,s6216,s6219);
  nand x3343(s6973,s6968,s6971);
  nand x3344(s7031,s7026,s7029);
  not x3345(s5521,s5515);
  nand x3346(s1756,s5515,s5522);
  not x3347(s5579,s5573);
  nand x3348(s1761,s5573,s5580);
  nand x3349(s5071,s5069,s5070);
  nand x3350(s5159,s5157,s5158);
  nand x3351(s5641,s5639,s5640);
  nand x3352(s5729,s5727,s5728);
  nand x3353(s6107,s6105,s6106);
  nand x3354(s6165,s6163,s6164);
  nand x3355(s6223,s6221,s6222);
  not x3356(s6317,s6311);
  nand x3357(s6320,s6311,s6318);
  nand x3358(s6975,s6973,s6974);
  nand x3359(s7033,s7031,s7032);
  not x3360(s7097,s7091);
  nand x3361(s7100,s7091,s7098);
  not x3362(s7185,s7179);
  nand x3363(s7188,s7179,s7186);
  nand x3364(s1755,s5518,s5521);
  nand x3365(s1760,s5576,s5579);
  nand x3366(s6319,s6314,s6317);
  nand x3367(s7099,s7094,s7097);
  nand x3368(s7187,s7182,s7185);
  nand x3369(s1757,s1755,s1756);
  nand x3370(s1762,s1760,s1761);
  not x3371(s6113,s6107);
  nand x3372(s2818,s6107,s6114);
  not x3373(s6171,s6165);
  nand x3374(s2823,s6165,s6172);
  not x3375(s6981,s6975);
  nand x3376(s4058,s6975,s6982);
  not x3377(s7039,s7033);
  nand x3378(s4063,s7033,s7040);
  not x3379(s5077,s5071);
  nand x3380(s5080,s5071,s5078);
  not x3381(s5165,s5159);
  nand x3382(s5090,s5159,s5166);
  not x3383(s5647,s5641);
  nand x3384(s5650,s5641,s5648);
  not x3385(s5735,s5729);
  nand x3386(s5660,s5729,s5736);
  not x3387(s6229,s6223);
  nand x3388(s6232,s6223,s6230);
  nand x3389(s6321,s6319,s6320);
  nand x3390(s7101,s7099,s7100);
  nand x3391(s7189,s7187,s7188);
  nand x3392(s2817,s6110,s6113);
  nand x3393(s2822,s6168,s6171);
  nand x3394(s4057,s6978,s6981);
  nand x3395(s4062,s7036,s7039);
  nand x3396(s5079,s5074,s5077);
  nand x3397(s5089,s5162,s5165);
  nand x3398(s5649,s5644,s5647);
  nand x3399(s5659,s5732,s5735);
  nand x3400(s6231,s6226,s6229);
  and x3401(s1782,s1762,s1730,s1771);
  and x3402(s1783,s1757,s1726,s1771);
  and x3403(s1784,s1762,s1751,s1766);
  and x3404(s1785,s1757,s1754,s1766);
  nand x3405(s2819,s2817,s2818);
  nand x3406(s2824,s2822,s2823);
  nand x3407(s4059,s4057,s4058);
  nand x3408(s4064,s4062,s4063);
  nand x3409(s5081,s5079,s5080);
  nand x3410(s5091,s5089,s5090);
  nand x3411(s5651,s5649,s5650);
  nand x3412(s5661,s5659,s5660);
  nand x3413(s6233,s6231,s6232);
  not x3414(s6327,s6321);
  nand x3415(s6252,s6321,s6328);
  not x3416(s7107,s7101);
  nand x3417(s7110,s7101,s7108);
  not x3418(s7195,s7189);
  nand x3419(s7120,s7189,s7196);
  or x3420(s5737,s1782,s1783,s1784,s1785);
  nand x3421(s6251,s6324,s6327);
  nand x3422(s7109,s7104,s7107);
  nand x3423(s7119,s7192,s7195);
  not x3424(s5087,s5081);
  nand x3425(s985,s5081,s5088);
  not x3426(s5097,s5091);
  nand x3427(s988,s5091,s5098);
  not x3428(s5657,s5651);
  nand x3429(s1776,s5651,s5658);
  not x3430(s5667,s5661);
  nand x3431(s1779,s5661,s5668);
  and x3432(s2844,s2824,s2784,s2833);
  and x3433(s2845,s2819,s2780,s2833);
  and x3434(s2846,s2824,s2813,s2828);
  and x3435(s2847,s2819,s2816,s2828);
  and x3436(s4083,s4064,s4032,s4072);
  and x3437(s4084,s4059,s4028,s4072);
  and x3438(s4085,s4064,s4053,s4067);
  and x3439(s4086,s4059,s4056,s4067);
  not x3440(s6239,s6233);
  nand x3441(s6242,s6233,s6240);
  nand x3442(s6253,s6251,s6252);
  nand x3443(s7111,s7109,s7110);
  nand x3444(s7121,s7119,s7120);
  nand x3445(s984,s5084,s5087);
  nand x3446(s987,s5094,s5097);
  nand x3447(s1775,s5654,s5657);
  nand x3448(s1778,s5664,s5667);
  not x3449(s5743,s5737);
  nand x3450(s6241,s6236,s6239);
  or x3451(s6329,s2844,s2845,s2846,s2847);
  or x3452(s7197,s4083,s4084,s4085,s4086);
  nand x3453(s986,s984,s985);
  nand x3454(s989,s987,s988);
  nand x3455(s1777,s1775,s1776);
  nand x3456(s1780,s1778,s1779);
  not x3457(s6259,s6253);
  nand x3458(s2841,s6253,s6260);
  not x3459(s7117,s7111);
  nand x3460(s4077,s7111,s7118);
  not x3461(s7127,s7121);
  nand x3462(s4080,s7121,s7128);
  nand x3463(s6243,s6241,s6242);
  not x3464(s990,s989);
  and x3465(s996,s975,s986);
  not x3466(s1781,s1780);
  and x3467(s1787,s1766,s1777);
  nand x3468(s2840,s6256,s6259);
  not x3469(s6335,s6329);
  nand x3470(s4076,s7114,s7117);
  nand x3471(s4079,s7124,s7127);
  not x3472(s7203,s7197);
  and x3473(s995,s990,s980);
  and x3474(s1786,s1781,s1771);
  not x3475(s6249,s6243);
  nand x3476(s2838,s6243,s6250);
  nand x3477(s2842,s2840,s2841);
  nand x3478(s4078,s4076,s4077);
  nand x3479(s4081,s4079,s4080);
  nand x3480(s2837,s6246,s6249);
  not x3481(s2843,s2842);
  not x3482(s4082,s4081);
  and x3483(s4088,s4067,s4078);
  or x3484(s5170,s995,s996);
  or x3485(s5740,s1786,s1787);
  nand x3486(s2839,s2837,s2838);
  and x3487(s2848,s2843,s2833);
  and x3488(s4087,s4082,s4072);
  nand x3489(s1791,s5740,s5743);
  nand x3490(s1003,s5170,s5173);
  not x3491(s5174,s5170);
  not x3492(s5744,s5740);
  and x3493(s2849,s2828,s2839);
  or x3494(s7200,s4087,s4088);
  nand x3495(s1792,s5737,s5744);
  nand x3496(s1004,s5167,s5174);
  or x3497(s6332,s2848,s2849);
  nand x3498(s320,s1791,s1792);
  nand x3499(s337,s1003,s1004);
  nand x3500(s4092,s7200,s7203);
  not x3501(s7204,s7200);
  not x3502(s321,s320);
  not x3503(s338,s337);
  nand x3504(s4093,s7197,s7204);
  nand x3505(s2855,s6332,s6335);
  not x3506(s6336,s6332);
  nand x3507(s369,s4092,s4093);
  nand x3508(s2856,s6329,s6336);
  not x3509(s370,s369);
  nand x3510(s398,s2855,s2856);
  not x3511(s399,s398);

endmodule
