module c1908(s3,s6,s9,s12,s30,s45,s48,s15,s18,s21,s24,s27,s33,s36,s39,s42,s75,s51,s54,s60,s63,s66,s69,s72,s57,s101,s104,s107,s110,s113,s116,s119,s122,s125,s128,s131,s134,s137,s140,s143,s146,s210,s214,s217,s221,s224,s227,s234,s237,s469,s472,s475,s478,s898,s900,s902,s952,s953);

  output s3;
  output s6;
  output s9;
  output s12;
  output s30;
  output s45;
  output s48;
  output s15;
  output s18;
  output s21;
  output s24;
  output s27;
  output s33;
  output s36;
  output s39;
  output s42;
  output s75;
  output s51;
  output s54;
  output s60;
  output s63;
  output s66;
  output s69;
  output s72;
  output s57;
  input s101;
  input s104;
  input s107;
  input s110;
  input s113;
  input s116;
  input s119;
  input s122;
  input s125;
  input s128;
  input s131;
  input s134;
  input s137;
  input s140;
  input s143;
  input s146;
  input s210;
  input s214;
  input s217;
  input s221;
  input s224;
  input s227;
  input s234;
  input s237;
  input s469;
  input s472;
  input s475;
  input s478;
  input s898;
  input s900;
  input s902;
  input s952;
  input s953;

  not x0(s149,s101);
  not x1(s153,s104);
  not x2(s156,s107);
  not x3(s160,s110);
  not x4(s165,s113);
  not x5(s168,s116);
  not x6(s171,s119);
  not x7(s175,s122);
  not x8(s179,s125);
  not x9(s184,s128);
  not x10(s188,s131);
  not x11(s191,s134);
  not x12(s194,s137);
  not x13(s198,s140);
  not x14(s202,s143);
  not x15(s206,s146);
  nand x16(s231,s224,s898);
  nand x17(s233,s227,s900);
  not x18(s241,s237);
  not x19(s244,s237);
  buf x20(s245,s234);
  buf x21(s248,s234);
  not x22(s517,s469);
  not x23(s529,s472);
  not x24(s541,s475);
  not x25(s553,s478);
  not x26(s859,s953);
  not x27(s862,s953);
  not x28(s907,s898);
  not x29(s909,s900);
  buf x30(s911,s902);
  not x31(s918,s902);
  buf x32(s919,s902);
  not x33(s922,s902);
  buf x34(s926,s952);
  not x35(s930,s952);
  not x36(s932,s952);
  buf x37(s934,s953);
  not x38(s938,s953);
  buf x39(s943,s953);
  buf x40(s947,s953);
  not x41(s949,s953);
  buf x42(s1506,s101);
  buf x43(s1514,s104);
  buf x44(s1522,s107);
  buf x45(s1530,s110);
  buf x46(s1538,s113);
  buf x47(s1546,s116);
  buf x48(s1554,s119);
  buf x49(s1562,s122);
  buf x50(s1570,s125);
  buf x51(s1578,s128);
  buf x52(s1586,s131);
  buf x53(s1594,s134);
  buf x54(s1602,s137);
  buf x55(s1610,s140);
  buf x56(s1618,s143);
  buf x57(s1626,s146);
  not x58(s1512,s1506);
  not x59(s1520,s1514);
  not x60(s1528,s1522);
  not x61(s1536,s1530);
  not x62(s1544,s1538);
  not x63(s1552,s1546);
  not x64(s1560,s1554);
  not x65(s1568,s1562);
  not x66(s1576,s1570);
  not x67(s1584,s1578);
  not x68(s1592,s1586);
  not x69(s1600,s1594);
  not x70(s1608,s1602);
  not x71(s1616,s1610);
  not x72(s1624,s1618);
  not x73(s1632,s1626);
  nand x74(s50,s930,s947);
  nand x75(s52,s930,s947);
  nand x76(s56,s930,s947);
  nand x77(s58,s930,s947);
  nand x78(s62,s930,s947);
  nand x79(s64,s930,s947);
  buf x80(s251,s149);
  buf x81(s254,s153);
  buf x82(s288,s165);
  buf x83(s291,s168);
  buf x84(s299,s184);
  buf x85(s302,s202);
  and x86(s318,s224,s938);
  buf x87(s321,s179);
  buf x88(s327,s188);
  buf x89(s330,s191);
  and x90(s352,s227,s938);
  buf x91(s355,s198);
  and x92(s369,s210,s241,s938);
  buf x93(s382,s206);
  buf x94(s385,s198);
  nand x95(s853,s943,s907);
  nand x96(s856,s943,s909);
  nand x97(s893,s248,s237);
  nand x98(s954,s248,s922);
  nand x99(s955,s244,s922);
  buf x100(s1050,s160);
  buf x101(s1053,s175);
  buf x102(s1176,s179);
  buf x103(s1179,s198);
  buf x104(s1197,s149);
  buf x105(s1207,s149);
  buf x106(s1222,s153);
  buf x107(s1244,s188);
  buf x108(s1278,s156);
  and x109(s1290,s217,s245,s938);
  buf x110(s1300,s191);
  buf x111(s1312,s160);
  buf x112(s1332,s194);
  and x113(s1335,s221,s245,s938);
  buf x114(s1442,s517);
  buf x115(s1450,s517);
  buf x116(s1458,s529);
  buf x117(s1466,s529);
  buf x118(s1474,s541);
  buf x119(s1482,s541);
  buf x120(s1490,s553);
  buf x121(s1498,s553);
  and x122(s1634,s231,s934);
  and x123(s1644,s233,s934);
  buf x124(s1657,s156);
  buf x125(s1665,s156);
  buf x126(s1697,s171);
  buf x127(s1705,s171);
  buf x128(s1713,s206);
  buf x129(s1721,s206);
  buf x130(s1745,s194);
  buf x131(s1753,s194);
  buf x132(s1785,s160);
  buf x133(s1793,s160);
  buf x134(s1814,s165);
  buf x135(s1817,s175);
  and x136(s1830,s214,s241,s938);
  buf x137(s1833,s202);
  buf x138(s1841,s179);
  buf x139(s1849,s179);
  buf x140(s1854,s168);
  buf x141(s1857,s175);
  buf x142(s1870,s184);
  buf x143(s1873,s202);
  buf x144(s1878,s171);
  buf x145(s1881,s184);
  not x146(s1642,s1634);
  not x147(s1652,s1644);
  not x148(s1056,s1050);
  not x149(s1057,s1053);
  not x150(s1182,s1176);
  not x151(s1183,s1179);
  not x152(s1211,s1207);
  not x153(s1298,s1290);
  not x154(s1320,s1312);
  not x155(s1338,s1332);
  not x156(s1339,s1335);
  and x157(s457,s210,s955);
  and x158(s459,s217,s954);
  nand x159(s482,s214,s955);
  nand x160(s487,s221,s954);
  nand x161(s492,s210,s955);
  nand x162(s505,s217,s954);
  not x163(s1456,s1450);
  not x164(s1448,s1442);
  not x165(s1472,s1466);
  not x166(s1464,s1458);
  not x167(s1488,s1482);
  not x168(s1480,s1474);
  not x169(s1504,s1498);
  not x170(s1496,s1490);
  nand x171(s956,s907,s919,s943,s893);
  nand x172(s967,s909,s919,s943,s893);
  nand x173(s978,s926,s949,s893);
  and x174(s979,s926,s949,s893);
  buf x175(s980,s251);
  not x176(s1661,s1657);
  buf x177(s990,s251);
  not x178(s1669,s1665);
  buf x179(s1030,s288);
  not x180(s1701,s1697);
  buf x181(s1040,s288);
  not x182(s1709,s1705);
  buf x183(s1058,s299);
  not x184(s1717,s1713);
  buf x185(s1068,s299);
  not x186(s1725,s1721);
  buf x187(s1078,s318);
  buf x188(s1090,s318);
  buf x189(s1100,s327);
  not x190(s1749,s1745);
  buf x191(s1112,s327);
  not x192(s1757,s1753);
  buf x193(s1154,s352);
  not x194(s1789,s1785);
  buf x195(s1166,s352);
  not x196(s1797,s1793);
  buf x197(s1194,s369);
  not x198(s1201,s1197);
  buf x199(s1204,s369);
  not x200(s1820,s1814);
  not x201(s1821,s1817);
  not x202(s1230,s1222);
  not x203(s1836,s1830);
  not x204(s1837,s1833);
  not x205(s1252,s1244);
  buf x206(s1256,s382);
  not x207(s1845,s1841);
  buf x208(s1268,s382);
  not x209(s1853,s1849);
  not x210(s1860,s1854);
  not x211(s1861,s1857);
  not x212(s1286,s1278);
  not x213(s1876,s1870);
  not x214(s1877,s1873);
  not x215(s1308,s1300);
  not x216(s1884,s1878);
  not x217(s1885,s1881);
  buf x218(s1654,s254);
  buf x219(s1662,s254);
  buf x220(s1694,s291);
  buf x221(s1702,s291);
  buf x222(s1710,s302);
  buf x223(s1718,s302);
  buf x224(s1726,s321);
  buf x225(s1734,s321);
  buf x226(s1742,s330);
  buf x227(s1750,s330);
  buf x228(s1782,s355);
  buf x229(s1790,s355);
  buf x230(s1838,s385);
  buf x231(s1846,s385);
  nand x232(s297,s1053,s1056);
  nand x233(s298,s1050,s1057);
  nand x234(s361,s1179,s1182);
  nand x235(s362,s1176,s1183);
  nand x236(s404,s1335,s1338);
  nand x237(s405,s1332,s1339);
  nand x238(s1225,s1817,s1820);
  nand x239(s1226,s1814,s1821);
  nand x240(s1247,s1833,s1836);
  nand x241(s1248,s1830,s1837);
  nand x242(s1281,s1857,s1860);
  nand x243(s1282,s1854,s1861);
  nand x244(s1303,s1873,s1876);
  nand x245(s1304,s1870,s1877);
  nand x246(s1315,s1881,s1884);
  nand x247(s1316,s1878,s1885);
  not x248(s998,s990);
  not x249(s988,s980);
  nand x250(s268,s297,s298);
  not x251(s1038,s1030);
  not x252(s1048,s1040);
  not x253(s1076,s1068);
  not x254(s1066,s1058);
  not x255(s1098,s1090);
  not x256(s1120,s1112);
  not x257(s1174,s1166);
  nand x258(s363,s361,s362);
  not x259(s1210,s1204);
  nand x260(s373,s1204,s1211);
  not x261(s1276,s1268);
  nand x262(s406,s404,s405);
  not x263(s565,s482);
  buf x264(s566,s482);
  not x265(s614,s487);
  buf x266(s615,s487);
  nand x267(s958,s956,s978);
  nand x268(s969,s967,s978);
  not x269(s1660,s1654);
  nand x270(s984,s1654,s1661);
  not x271(s1668,s1662);
  nand x272(s994,s1662,s1669);
  not x273(s1700,s1694);
  nand x274(s1034,s1694,s1701);
  not x275(s1708,s1702);
  nand x276(s1044,s1702,s1709);
  not x277(s1716,s1710);
  nand x278(s1062,s1710,s1717);
  not x279(s1724,s1718);
  nand x280(s1072,s1718,s1725);
  not x281(s1732,s1726);
  not x282(s1086,s1078);
  not x283(s1740,s1734);
  not x284(s1748,s1742);
  nand x285(s1104,s1742,s1749);
  not x286(s1108,s1100);
  not x287(s1756,s1750);
  nand x288(s1116,s1750,s1757);
  not x289(s1788,s1782);
  nand x290(s1158,s1782,s1789);
  not x291(s1162,s1154);
  not x292(s1796,s1790);
  nand x293(s1170,s1790,s1797);
  not x294(s1200,s1194);
  nand x295(s1203,s1194,s1201);
  nand x296(s1227,s1225,s1226);
  nand x297(s1249,s1247,s1248);
  not x298(s1844,s1838);
  nand x299(s1260,s1838,s1845);
  not x300(s1264,s1256);
  not x301(s1852,s1846);
  nand x302(s1272,s1846,s1853);
  nand x303(s1283,s1281,s1282);
  nand x304(s1305,s1303,s1304);
  nand x305(s1317,s1315,s1316);
  buf x306(s1410,s492);
  buf x307(s1418,s492);
  buf x308(s1426,s505);
  buf x309(s1434,s505);
  not x310(s269,s268);
  nand x311(s372,s1207,s1210);
  nand x312(s983,s1657,s1660);
  nand x313(s993,s1665,s1668);
  nand x314(s1033,s1697,s1700);
  nand x315(s1043,s1705,s1708);
  nand x316(s1061,s1713,s1716);
  nand x317(s1071,s1721,s1724);
  nand x318(s1103,s1745,s1748);
  nand x319(s1115,s1753,s1756);
  nand x320(s1157,s1785,s1788);
  nand x321(s1169,s1793,s1796);
  not x322(s1184,s363);
  nand x323(s1202,s1197,s1200);
  nand x324(s1259,s1841,s1844);
  nand x325(s1271,s1849,s1852);
  not x326(s1322,s406);
  nand x327(s374,s372,s373);
  nand x328(s396,s1317,s1320);
  not x329(s1321,s1317);
  not x330(s1424,s1418);
  not x331(s1416,s1410);
  not x332(s1440,s1434);
  not x333(s1432,s1426);
  nand x334(s985,s983,s984);
  nand x335(s995,s993,s994);
  nand x336(s1035,s1033,s1034);
  nand x337(s1045,s1043,s1044);
  nand x338(s1063,s1061,s1062);
  nand x339(s1073,s1071,s1072);
  nand x340(s1105,s1103,s1104);
  nand x341(s1117,s1115,s1116);
  nand x342(s1159,s1157,s1158);
  nand x343(s1171,s1169,s1170);
  nand x344(s1212,s1202,s1203);
  not x345(s1231,s1227);
  nand x346(s1232,s1227,s1230);
  not x347(s1253,s1249);
  nand x348(s1254,s1249,s1252);
  nand x349(s1261,s1259,s1260);
  nand x350(s1273,s1271,s1272);
  not x351(s1287,s1283);
  nand x352(s1288,s1283,s1286);
  not x353(s1309,s1305);
  nand x354(s1310,s1305,s1308);
  not x355(s1192,s1184);
  nand x356(s397,s1312,s1321);
  not x357(s1330,s1322);
  buf x358(s1000,s269);
  buf x359(s1010,s269);
  nand x360(s1233,s1222,s1231);
  nand x361(s1255,s1244,s1253);
  nand x362(s1289,s1278,s1287);
  nand x363(s1311,s1300,s1309);
  not x364(s1381,s374);
  nand x365(s257,s995,s998);
  not x366(s999,s995);
  nand x367(s260,s985,s988);
  not x368(s989,s985);
  nand x369(s272,s1035,s1038);
  not x370(s1039,s1035);
  nand x371(s294,s1045,s1048);
  not x372(s1049,s1045);
  nand x373(s305,s1073,s1076);
  not x374(s1077,s1073);
  nand x375(s308,s1063,s1066);
  not x376(s1067,s1063);
  nand x377(s333,s1117,s1120);
  not x378(s1121,s1117);
  nand x379(s358,s1171,s1174);
  not x380(s1175,s1171);
  not x381(s1220,s1212);
  nand x382(s388,s1273,s1276);
  not x383(s1277,s1273);
  nand x384(s398,s396,s397);
  not x385(s1109,s1105);
  nand x386(s1110,s1105,s1108);
  not x387(s1163,s1159);
  nand x388(s1164,s1159,s1162);
  nand x389(s1234,s1232,s1233);
  not x390(s1265,s1261);
  nand x391(s1266,s1261,s1264);
  nand x392(s1822,s1254,s1255);
  nand x393(s1862,s1310,s1311);
  nand x394(s1865,s1288,s1289);
  nand x395(s258,s990,s999);
  nand x396(s261,s980,s989);
  nand x397(s273,s1030,s1039);
  not x398(s1018,s1010);
  not x399(s1008,s1000);
  nand x400(s295,s1040,s1049);
  nand x401(s306,s1068,s1077);
  nand x402(s309,s1058,s1067);
  nand x403(s334,s1112,s1121);
  nand x404(s359,s1166,s1175);
  nand x405(s389,s1268,s1277);
  not x406(s1385,s1381);
  nand x407(s1111,s1100,s1109);
  nand x408(s1165,s1154,s1163);
  nand x409(s1267,s1256,s1265);
  not x410(s1886,s398);
  nand x411(s259,s257,s258);
  nand x412(s262,s260,s261);
  nand x413(s274,s272,s273);
  nand x414(s296,s294,s295);
  nand x415(s307,s305,s306);
  nand x416(s310,s308,s309);
  nand x417(s335,s333,s334);
  nand x418(s360,s358,s359);
  not x419(s1242,s1234);
  nand x420(s390,s388,s389);
  not x421(s1828,s1822);
  not x422(s1868,s1862);
  not x423(s1869,s1865);
  nand x424(s1373,s1164,s1165);
  nand x425(s1798,s1110,s1111);
  nand x426(s1825,s1266,s1267);
  not x427(s265,s259);
  not x428(s314,s307);
  not x429(s336,s335);
  not x430(s407,s296);
  nand x431(s1293,s1865,s1868);
  nand x432(s1294,s1862,s1869);
  not x433(s1892,s1886);
  not x434(s1777,s360);
  not x435(s1889,s390);
  buf x436(s410,s310);
  not x437(s1377,s1373);
  not x438(s1804,s1798);
  nand x439(s1237,s1825,s1828);
  not x440(s1829,s1825);
  nand x441(s1295,s1293,s1294);
  buf x442(s1670,s274);
  buf x443(s1678,s274);
  buf x444(s1729,s310);
  buf x445(s1737,s310);
  buf x446(s1761,s262);
  buf x447(s1769,s262);
  buf x448(s340,s336);
  buf x449(s343,s314);
  not x450(s1781,s1777);
  nand x451(s1238,s1822,s1829);
  nand x452(s1325,s1889,s1892);
  not x453(s1893,s1889);
  buf x454(s1340,s407);
  buf x455(s1352,s407);
  buf x456(s1673,s265);
  buf x457(s1681,s265);
  buf x458(s1801,s314);
  buf x459(s1897,s336);
  buf x460(s1905,s336);
  nand x461(s391,s1295,s1298);
  not x462(s1299,s1295);
  not x463(s1676,s1670);
  not x464(s1684,s1678);
  nand x465(s1081,s1729,s1732);
  not x466(s1733,s1729);
  nand x467(s1093,s1737,s1740);
  not x468(s1741,s1737);
  not x469(s1765,s1761);
  not x470(s1773,s1769);
  nand x471(s1239,s1237,s1238);
  nand x472(s1326,s1886,s1893);
  buf x473(s1894,s410);
  buf x474(s1902,s410);
  nand x475(s392,s1290,s1299);
  not x476(s1360,s1352);
  nand x477(s1003,s1673,s1676);
  not x478(s1677,s1673);
  nand x479(s1013,s1681,s1684);
  not x480(s1685,s1681);
  nand x481(s1082,s1726,s1733);
  nand x482(s1094,s1734,s1741);
  buf x483(s1122,s340);
  buf x484(s1134,s340);
  nand x485(s1187,s1801,s1804);
  not x486(s1805,s1801);
  nand x487(s1327,s1325,s1326);
  not x488(s1901,s1897);
  not x489(s1348,s1340);
  not x490(s1909,s1905);
  buf x491(s1758,s343);
  buf x492(s1766,s343);
  nand x493(s377,s1239,s1242);
  not x494(s1243,s1239);
  nand x495(s393,s391,s392);
  nand x496(s1004,s1670,s1677);
  nand x497(s1014,s1678,s1685);
  nand x498(s1083,s1081,s1082);
  nand x499(s1095,s1093,s1094);
  nand x500(s1188,s1798,s1805);
  not x501(s1900,s1894);
  nand x502(s1344,s1894,s1901);
  not x503(s1908,s1902);
  nand x504(s1356,s1902,s1909);
  not x505(s1142,s1134);
  nand x506(s378,s1234,s1243);
  nand x507(s399,s1327,s1330);
  not x508(s1331,s1327);
  nand x509(s1005,s1003,s1004);
  nand x510(s1015,s1013,s1014);
  not x511(s1764,s1758);
  nand x512(s1126,s1758,s1765);
  not x513(s1130,s1122);
  not x514(s1772,s1766);
  nand x515(s1138,s1766,s1773);
  nand x516(s1189,s1187,s1188);
  nand x517(s1343,s1897,s1900);
  nand x518(s1355,s1905,s1908);
  nand x519(s324,s1095,s1098);
  not x520(s1099,s1095);
  nand x521(s379,s377,s378);
  nand x522(s400,s1322,s1331);
  nand x523(s449,s393,s918);
  not x524(s1087,s1083);
  nand x525(s1088,s1083,s1086);
  nand x526(s1125,s1761,s1764);
  nand x527(s1137,s1769,s1772);
  nand x528(s1345,s1343,s1344);
  nand x529(s1357,s1355,s1356);
  buf x530(s1397,s393);
  nand x531(s277,s1015,s1018);
  not x532(s1019,s1015);
  nand x533(s280,s1005,s1008);
  not x534(s1009,s1005);
  nand x535(s325,s1090,s1099);
  nand x536(s364,s1189,s1192);
  not x537(s1193,s1189);
  nand x538(s401,s399,s400);
  nand x539(s1089,s1078,s1087);
  nand x540(s1127,s1125,s1126);
  nand x541(s1139,s1137,s1138);
  nand x542(s278,s1010,s1019);
  nand x543(s281,s1000,s1009);
  nand x544(s326,s324,s325);
  nand x545(s365,s1184,s1193);
  nand x546(s413,s1357,s1360);
  not x547(s1361,s1357);
  not x548(s1401,s1397);
  nand x549(s445,s379,s918);
  not x550(s1349,s1345);
  nand x551(s1350,s1345,s1348);
  buf x552(s1389,s379);
  buf x553(s1493,s449);
  buf x554(s1501,s449);
  nand x555(s1689,s1088,s1089);
  nand x556(s279,s277,s278);
  nand x557(s282,s280,s281);
  nand x558(s346,s1139,s1142);
  not x559(s1143,s1139);
  nand x560(s366,s364,s365);
  nand x561(s414,s1352,s1361);
  nand x562(s453,s401,s918);
  not x563(s1131,s1127);
  nand x564(s1132,s1127,s1130);
  nand x565(s1351,s1340,s1349);
  not x566(s1365,s326);
  buf x567(s1405,s401);
  not x568(s285,s279);
  nand x569(s347,s1134,s1143);
  not x570(s367,s366);
  nand x571(s415,s413,s414);
  not x572(s1393,s1389);
  nand x573(s556,s1501,s1504);
  not x574(s1505,s1501);
  nand x575(s559,s1493,s1496);
  not x576(s1497,s1493);
  not x577(s1693,s1689);
  nand x578(s1133,s1122,s1131);
  buf x579(s1477,s445);
  buf x580(s1485,s445);
  nand x581(s1809,s1350,s1351);
  nand x582(s348,s346,s347);
  not x583(s1369,s1365);
  not x584(s1409,s1405);
  nand x585(s557,s1498,s1505);
  nand x586(s560,s1490,s1497);
  buf x587(s1362,s282);
  not x588(s1378,s415);
  buf x589(s1429,s453);
  buf x590(s1437,s453);
  buf x591(s1686,s282);
  nand x592(s1774,s1132,s1133);
  and x593(s1910,s285,s853);
  and x594(s1918,s856,s367);
  nand x595(s544,s1485,s1488);
  not x596(s1489,s1485);
  nand x597(s547,s1477,s1480);
  not x598(s1481,s1477);
  nand x599(s558,s556,s557);
  nand x600(s561,s559,s560);
  not x601(s1813,s1809);
  not x602(s1370,s348);
  not x603(s1368,s1362);
  nand x604(s417,s1362,s1369);
  not x605(s1384,s1378);
  nand x606(s424,s1378,s1385);
  nand x607(s508,s1437,s1440);
  not x608(s1441,s1437);
  nand x609(s511,s1429,s1432);
  not x610(s1433,s1429);
  nand x611(s545,s1482,s1489);
  nand x612(s548,s1474,s1481);
  not x613(s564,s558);
  not x614(s1692,s1686);
  nand x615(s1024,s1686,s1693);
  not x616(s1780,s1774);
  nand x617(s1148,s1774,s1781);
  not x618(s1916,s1910);
  not x619(s1924,s1918);
  nand x620(s416,s1365,s1368);
  not x621(s1376,s1370);
  nand x622(s421,s1370,s1377);
  nand x623(s423,s1381,s1384);
  nand x624(s509,s1434,s1441);
  nand x625(s512,s1426,s1433);
  nand x626(s546,s544,s545);
  nand x627(s549,s547,s548);
  not x628(s719,s561);
  buf x629(s722,s561);
  nand x630(s1023,s1689,s1692);
  nand x631(s1147,s1777,s1780);
  nand x632(s418,s416,s417);
  nand x633(s420,s1373,s1376);
  nand x634(s425,s423,s424);
  nand x635(s510,s508,s509);
  nand x636(s513,s511,s512);
  not x637(s552,s546);
  nand x638(s1025,s1023,s1024);
  nand x639(s1149,s1147,s1148);
  not x640(s419,s418);
  nand x641(s422,s420,s421);
  nand x642(s441,s425,s918);
  not x643(s516,s510);
  not x644(s725,s549);
  buf x645(s728,s549);
  not x646(s1029,s1025);
  not x647(s1153,s1149);
  nand x648(s433,s419,s918);
  nand x649(s437,s422,s918);
  not x650(s663,s513);
  buf x651(s666,s513);
  and x652(s731,s719,s725);
  and x653(s746,s722,s725);
  and x654(s756,s719,s728);
  and x655(s770,s722,s728);
  buf x656(s1461,s441);
  buf x657(s1469,s441);
  buf x658(s1413,s433);
  buf x659(s1421,s433);
  buf x660(s1445,s437);
  buf x661(s1453,s437);
  nand x662(s532,s1469,s1472);
  not x663(s1473,s1469);
  nand x664(s535,s1461,s1464);
  not x665(s1465,s1461);
  nand x666(s495,s1421,s1424);
  not x667(s1425,s1421);
  nand x668(s498,s1413,s1416);
  not x669(s1417,s1413);
  nand x670(s520,s1453,s1456);
  not x671(s1457,s1453);
  nand x672(s523,s1445,s1448);
  not x673(s1449,s1445);
  nand x674(s533,s1466,s1473);
  nand x675(s536,s1458,s1465);
  nand x676(s496,s1418,s1425);
  nand x677(s499,s1410,s1417);
  nand x678(s521,s1450,s1457);
  nand x679(s524,s1442,s1449);
  nand x680(s534,s532,s533);
  nand x681(s537,s535,s536);
  nand x682(s497,s495,s496);
  nand x683(s500,s498,s499);
  nand x684(s522,s520,s521);
  nand x685(s525,s523,s524);
  not x686(s540,s534);
  not x687(s503,s497);
  not x688(s528,s522);
  not x689(s669,s537);
  buf x690(s672,s537);
  not x691(s569,s500);
  and x692(s588,s566,s500);
  not x693(s618,s525);
  and x694(s639,s615,s525);
  nand x695(s867,s516,s564,s552,s540,s482,s528,s503,s487);
  buf x696(s588a,s588);
  buf x697(s588b,s588);
  buf x698(s639a,s639);
  buf x699(s639b,s639);
  and x700(s675,s663,s669);
  and x701(s688,s666,s669);
  and x702(s696,s663,s672);
  and x703(s710,s666,s672);
  and x704(s73,s949,s867,s932,s932);
  and x705(s572,s565,s569);
  and x706(s573,s566,s569);
  and x707(s621,s614,s618);
  and x708(s622,s615,s618);
  nand x709(s776,s588a,s639a,s696,s731,s958);
  nand x710(s780,s588a,s639a,s675,s756,s958);
  nand x711(s784,s588a,s639a,s675,s746,s958);
  nand x712(s788,s588a,s639a,s688,s731,s958);
  nand x713(s812,s588b,s639a,s710,s746,s969);
  nand x714(s832,s588b,s639b,s696,s770,s969);
  nand x715(s836,s588b,s639b,s710,s756,s969);
  and x716(s1509,s588a,s639a,s696,s731,s958);
  and x717(s1517,s588a,s639a,s675,s756,s958);
  and x718(s1525,s588a,s639a,s675,s746,s958);
  and x719(s1533,s588a,s639a,s688,s731,s958);
  and x720(s1581,s588b,s639a,s710,s746,s969);
  and x721(s1621,s588b,s639b,s696,s770,s969);
  and x722(s1629,s588b,s639b,s710,s756,s969);
  nand x723(s792,s588a,s622,s696,s756,s958);
  nand x724(s796,s588b,s622,s696,s746,s958);
  nand x725(s800,s588b,s622,s710,s731,s958);
  nand x726(s804,s588b,s622,s675,s770,s958);
  nand x727(s808,s588b,s622,s688,s756,s969);
  nand x728(s816,s573,s639b,s696,s756,s969);
  nand x729(s820,s573,s639b,s696,s746,s969);
  nand x730(s824,s573,s639b,s710,s731,s969);
  nand x731(s828,s573,s639b,s688,s756,s969);
  nand x732(s871,s588b,s622,s675,s731,s979);
  nand x733(s873,s573,s639b,s675,s731,s979);
  nand x734(s875,s573,s622,s696,s731,s979);
  nand x735(s877,s573,s622,s675,s756,s979);
  nand x736(s879,s573,s622,s675,s746,s979);
  nand x737(s881,s573,s622,s688,s731,s979);
  nand x738(s883,s573,s621,s675,s731,s979);
  nand x739(s885,s572,s622,s675,s731,s979);
  and x740(s1541,s588a,s622,s696,s756,s958);
  and x741(s1549,s588b,s622,s696,s746,s958);
  and x742(s1557,s588b,s622,s710,s731,s958);
  and x743(s1565,s588b,s622,s675,s770,s958);
  and x744(s1573,s588b,s622,s688,s756,s969);
  and x745(s1589,s573,s639b,s696,s756,s969);
  and x746(s1597,s573,s639b,s696,s746,s969);
  and x747(s1605,s573,s639b,s710,s731,s969);
  and x748(s1613,s573,s639b,s688,s756,s969);
  nand x749(s1,s1509,s1512);
  not x750(s1513,s1509);
  nand x751(s4,s1517,s1520);
  not x752(s1521,s1517);
  nand x753(s7,s1525,s1528);
  not x754(s1529,s1525);
  nand x755(s10,s1533,s1536);
  not x756(s1537,s1533);
  nand x757(s28,s1581,s1584);
  not x758(s1585,s1581);
  nand x759(s43,s1621,s1624);
  not x760(s1625,s1621);
  nand x761(s46,s1629,s1632);
  not x762(s1633,s1629);
  and x763(s886,s871,s873,s875,s877,s879,s881,s883,s885);
  nand x764(s2,s1506,s1513);
  nand x765(s5,s1514,s1521);
  nand x766(s8,s1522,s1529);
  nand x767(s11,s1530,s1537);
  nand x768(s13,s1541,s1544);
  not x769(s1545,s1541);
  nand x770(s16,s1549,s1552);
  not x771(s1553,s1549);
  nand x772(s19,s1557,s1560);
  not x773(s1561,s1557);
  nand x774(s22,s1565,s1568);
  not x775(s1569,s1565);
  nand x776(s25,s1573,s1576);
  not x777(s1577,s1573);
  nand x778(s29,s1578,s1585);
  nand x779(s31,s1589,s1592);
  not x780(s1593,s1589);
  nand x781(s34,s1597,s1600);
  not x782(s1601,s1597);
  nand x783(s37,s1605,s1608);
  not x784(s1609,s1605);
  nand x785(s40,s1613,s1616);
  not x786(s1617,s1613);
  nand x787(s44,s1618,s1625);
  nand x788(s47,s1626,s1633);
  nand x789(s857,s776,s780,s784,s788,s792,s796,s800,s804);
  nand x790(s860,s808,s812,s816,s820,s824,s828,s832,s836);
  and x791(s863,s776,s780,s784,s788,s792,s796,s800,s804);
  and x792(s865,s808,s812,s816,s820,s824,s828,s832,s836);
  nand x793(s3,s1,s2);
  nand x794(s6,s4,s5);
  nand x795(s9,s7,s8);
  nand x796(s12,s10,s11);
  nand x797(s14,s1538,s1545);
  nand x798(s17,s1546,s1553);
  nand x799(s20,s1554,s1561);
  nand x800(s23,s1562,s1569);
  nand x801(s26,s1570,s1577);
  nand x802(s30,s28,s29);
  nand x803(s32,s1586,s1593);
  nand x804(s35,s1594,s1601);
  nand x805(s38,s1602,s1609);
  nand x806(s41,s1610,s1617);
  nand x807(s45,s43,s44);
  nand x808(s48,s46,s47);
  and x809(s1913,s857,s859);
  and x810(s1921,s860,s862);
  nand x811(s15,s13,s14);
  nand x812(s18,s16,s17);
  nand x813(s21,s19,s20);
  nand x814(s24,s22,s23);
  nand x815(s27,s25,s26);
  nand x816(s33,s31,s32);
  nand x817(s36,s34,s35);
  nand x818(s39,s37,s38);
  nand x819(s42,s40,s41);
  and x820(s887,s863,s865,s886);
  nand x821(s462,s863,s865);
  and x822(s74,s949,s867,s952,s887);
  nand x823(s1637,s1913,s1916);
  not x824(s1917,s1913);
  nand x825(s1647,s1921,s1924);
  not x826(s1925,s1921);
  nor x827(s75,s73,s74);
  and x828(s1020,s457,s911,s462);
  and x829(s1144,s469,s911,s462);
  and x830(s1386,s475,s911,s462);
  and x831(s1394,s478,s911,s462);
  and x832(s1402,s459,s911,s462);
  nand x833(s1638,s1910,s1917);
  nand x834(s1648,s1918,s1925);
  and x835(s1806,s472,s911,s462);
  nand x836(s1639,s1637,s1638);
  nand x837(s1649,s1647,s1648);
  nand x838(s287,s1020,s1029);
  nand x839(s350,s1144,s1153);
  nand x840(s427,s1386,s1393);
  nand x841(s429,s1394,s1401);
  nand x842(s431,s1402,s1409);
  not x843(s1028,s1020);
  not x844(s1152,s1144);
  not x845(s1392,s1386);
  not x846(s1400,s1394);
  not x847(s1408,s1402);
  not x848(s1812,s1806);
  nand x849(s1216,s1806,s1813);
  nand x850(s286,s1025,s1028);
  nand x851(s349,s1149,s1152);
  nand x852(s426,s1389,s1392);
  nand x853(s428,s1397,s1400);
  nand x854(s430,s1405,s1408);
  nand x855(s67,s1639,s1642);
  not x856(s1643,s1639);
  nand x857(s70,s1649,s1652);
  not x858(s1653,s1649);
  nand x859(s1215,s1809,s1812);
  nand x860(s49,s286,s287);
  nand x861(s53,s349,s350);
  nand x862(s59,s426,s427);
  nand x863(s61,s428,s429);
  nand x864(s65,s430,s431);
  nand x865(s68,s1634,s1643);
  nand x866(s71,s1644,s1653);
  nand x867(s1217,s1215,s1216);
  and x868(s51,s49,s50);
  and x869(s54,s52,s53);
  and x870(s60,s58,s59);
  and x871(s63,s61,s62);
  and x872(s66,s64,s65);
  nand x873(s69,s67,s68);
  nand x874(s72,s70,s71);
  nand x875(s375,s1217,s1220);
  not x876(s1221,s1217);
  nand x877(s376,s1212,s1221);
  nand x878(s55,s375,s376);
  and x879(s57,s55,s56);

endmodule
