module c3540(s353,s355,s361,s358,s351,s372,s369,s399,s364,s396,s384,s367,s387,s393,s390,s378,s375,s381,s407,s409,s405,s402,s1,s13,s20,s33,s41,s45,s50,s58,s68,s77,s87,s97,s107,s116,s124,s125,s128,s132,s137,s143,s150,s159,s169,s179,s190,s200,s213,s222,s223,s226,s232,s238,s244,s250,s257,s264,s270,s274,s283,s294,s303,s311,s317,s322,s326,s329,s330,s343,s1698,s2897);

  output s353;
  output s355;
  output s361;
  output s358;
  output s351;
  output s372;
  output s369;
  output s399;
  output s364;
  output s396;
  output s384;
  output s367;
  output s387;
  output s393;
  output s390;
  output s378;
  output s375;
  output s381;
  output s407;
  output s409;
  output s405;
  output s402;
  input s1;
  input s13;
  input s20;
  input s33;
  input s41;
  input s45;
  input s50;
  input s58;
  input s68;
  input s77;
  input s87;
  input s97;
  input s107;
  input s116;
  input s124;
  input s125;
  input s128;
  input s132;
  input s137;
  input s143;
  input s150;
  input s159;
  input s169;
  input s179;
  input s190;
  input s200;
  input s213;
  input s222;
  input s223;
  input s226;
  input s232;
  input s238;
  input s244;
  input s250;
  input s257;
  input s264;
  input s270;
  input s274;
  input s283;
  input s294;
  input s303;
  input s311;
  input s317;
  input s322;
  input s326;
  input s329;
  input s330;
  input s343;
  input s1698;
  input s2897;

  buf x0(s432,s50);
  not x1(s442,s50);
  buf x2(s447,s58);
  not x3(s456,s58);
  buf x4(s460,s68);
  not x5(s463,s68);
  buf x6(s467,s68);
  buf x7(s476,s77);
  not x8(s479,s77);
  buf x9(s483,s77);
  buf x10(s492,s87);
  not x11(s501,s87);
  buf x12(s504,s97);
  not x13(s513,s97);
  buf x14(s517,s107);
  not x15(s526,s107);
  buf x16(s530,s116);
  not x17(s540,s116);
  or x18(s587,s257,s264);
  not x19(s704,s1);
  buf x20(s707,s1);
  not x21(s714,s1);
  buf x22(s717,s13);
  not x23(s724,s13);
  and x24(s731,s13,s20);
  not x25(s732,s20);
  buf x26(s736,s20);
  not x27(s741,s20);
  not x28(s758,s33);
  buf x29(s776,s33);
  not x30(s780,s33);
  and x31(s788,s33,s41);
  not x32(s791,s41);
  or x33(s798,s41,s45);
  buf x34(s799,s45);
  not x35(s802,s45);
  not x36(s826,s50);
  buf x37(s828,s58);
  not x38(s831,s58);
  buf x39(s833,s68);
  not x40(s836,s68);
  buf x41(s839,s87);
  not x42(s842,s87);
  buf x43(s845,s97);
  not x44(s848,s97);
  not x45(s851,s107);
  buf x46(s890,s1);
  buf x47(s898,s68);
  buf x48(s907,s107);
  not x49(s1032,s20);
  buf x50(s1035,s190);
  not x51(s1048,s200);
  and x52(s1049,s20,s200);
  nand x53(s1050,s20,s200);
  and x54(s1051,s20,s179);
  not x55(s1540,s20);
  or x56(s1699,s1698,s33);
  nand x57(s1826,s1,s13);
  nand x58(s1827,s1,s20,s33);
  not x59(s1828,s20);
  not x60(s2051,s33);
  buf x61(s2478,s179);
  not x62(s2865,s213);
  buf x63(s2868,s343);
  buf x64(s2931,s226);
  buf x65(s2934,s232);
  buf x66(s2939,s238);
  buf x67(s2942,s244);
  buf x68(s2947,s250);
  buf x69(s2950,s257);
  buf x70(s2957,s264);
  buf x71(s2960,s270);
  buf x72(s3007,s50);
  buf x73(s3079,s58);
  buf x74(s3087,s58);
  buf x75(s3095,s97);
  buf x76(s3103,s97);
  buf x77(s3419,s330);
  and x78(s588,s250,s587);
  or x79(s759,s758,s20);
  or x80(s1541,s1540,s169);
  not x81(s1772,s731);
  or x82(s1829,s1828,s1);
  and x83(s1834,s1826,s1827);
  or x84(s2052,s2051,s1);
  and x85(s625,s826,s831,s836);
  nand x86(s545,s226,s432);
  nand x87(s546,s232,s447);
  nand x88(s547,s238,s467);
  nand x89(s548,s244,s483);
  nand x90(s549,s250,s492);
  nand x91(s550,s257,s504);
  nand x92(s551,s264,s517);
  nand x93(s552,s270,s530);
  not x94(s2937,s2931);
  not x95(s2938,s2934);
  not x96(s2945,s2939);
  not x97(s2946,s2942);
  nand x98(s621,s456,s463);
  nand x99(s626,s513,s526);
  nand x100(s635,s460,s476);
  buf x101(s636,s442);
  not x102(s3085,s3079);
  not x103(s3101,s3095);
  buf x104(s657,s802);
  buf x105(s675,s802);
  buf x106(s721,s717);
  buf x107(s784,s780);
  buf x108(s794,s791);
  and x109(s807,s714,s798);
  and x110(s816,s714,s799,s791);
  and x111(s823,s704,s799);
  and x112(s860,s707,s724,s736);
  nand x113(s861,s707,s724,s736);
  nand x114(s864,s707,s724);
  buf x115(s893,s890);
  nand x116(s896,s717,s732,s45);
  nand x117(s897,s826,s831,s836);
  not x118(s3093,s3087);
  and x119(s905,s842,s848,s851);
  nand x120(s906,s842,s848,s851);
  not x121(s3109,s3103);
  not x122(s973,s741);
  not x123(s980,s741);
  not x124(s987,s741);
  not x125(s994,s741);
  not x126(s1001,s741);
  not x127(s1008,s741);
  not x128(s1015,s741);
  not x129(s1022,s741);
  or x130(s1038,s1032,s1035);
  nor x131(s1043,s1032,s1035);
  buf x132(s1054,s1051);
  not x133(s1057,s1051);
  buf x134(s1512,s776);
  buf x135(s1681,s780);
  not x136(s1717,s1699);
  not x137(s1724,s1699);
  not x138(s1731,s1699);
  not x139(s1738,s1699);
  not x140(s1745,s1699);
  not x141(s1752,s1699);
  not x142(s1759,s1699);
  not x143(s1766,s1699);
  or x144(s1773,s1,s1772);
  not x145(s1790,s788);
  not x146(s1808,s788);
  and x147(s2278,s704,s717,s732);
  not x148(s2481,s2478);
  not x149(s3425,s3419);
  or x150(s2871,s2865,s2868);
  nor x151(s2874,s2865,s2868);
  not x152(s2953,s2947);
  not x153(s2954,s2950);
  not x154(s2963,s2957);
  not x155(s2964,s2960);
  buf x156(s3010,s456);
  not x157(s3013,s3007);
  buf x158(s3017,s463);
  buf x159(s3020,s479);
  buf x160(s3027,s501);
  buf x161(s3030,s513);
  buf x162(s3037,s526);
  buf x163(s3040,s540);
  buf x164(s3082,s898);
  buf x165(s3090,s898);
  buf x166(s3098,s907);
  buf x167(s3106,s907);
  nand x168(s352,s479,s625);
  and x169(s553,s545,s546,s547,s548);
  and x170(s554,s549,s550,s551,s552);
  nand x171(s555,s2934,s2937);
  nand x172(s556,s2931,s2938);
  nand x173(s560,s2942,s2945);
  nand x174(s561,s2939,s2946);
  and x175(s650,s432,s621);
  and x176(s956,s890,s896);
  not x177(s974,s759);
  and x178(s975,s741,s759);
  and x179(s976,s897,s973);
  not x180(s981,s759);
  and x181(s982,s741,s759);
  not x182(s988,s759);
  and x183(s989,s741,s759);
  and x184(s990,s836,s987);
  not x185(s995,s759);
  and x186(s996,s741,s759);
  and x187(s997,s77,s994);
  not x188(s1002,s759);
  and x189(s1003,s741,s759);
  and x190(s1004,s906,s1001);
  not x191(s1009,s759);
  and x192(s1010,s741,s759);
  not x193(s1016,s759);
  and x194(s1017,s741,s759);
  and x195(s1018,s851,s1015);
  not x196(s1023,s759);
  and x197(s1024,s741,s759);
  and x198(s1025,s116,s1022);
  and x199(s1720,s222,s1717);
  and x200(s1727,s223,s1724);
  and x201(s1734,s226,s1731);
  and x202(s1741,s232,s1738);
  and x203(s1748,s238,s1745);
  and x204(s1755,s244,s1752);
  and x205(s1762,s250,s1759);
  and x206(s1769,s257,s1766);
  and x207(s1791,s1,s13,s1790);
  and x208(s1809,s1,s13,s1808);
  not x209(s1851,s1834);
  not x210(s1901,s1834);
  not x211(s1952,s1834);
  not x212(s2002,s1834);
  not x213(s2057,s1834);
  not x214(s2109,s1834);
  not x215(s2162,s1834);
  not x216(s2214,s1834);
  nand x217(s2955,s2950,s2953);
  nand x218(s2956,s2947,s2954);
  nand x219(s2965,s2960,s2963);
  nand x220(s2966,s2957,s2964);
  not x221(s353,s352);
  and x222(s354,s87,s626);
  nand x223(s557,s555,s556);
  nand x224(s562,s560,s561);
  nand x225(s586,s553,s554);
  and x226(s630,s540,s905);
  nand x227(s634,s540,s905);
  not x228(s639,s636);
  nand x229(s642,s3082,s3085);
  not x230(s3086,s3082);
  and x231(s644,s460,s636);
  nand x232(s646,s3098,s3101);
  not x233(s3102,s3098);
  nand x234(s654,s87,s626);
  not x235(s660,s657);
  not x236(s678,s675);
  nand x237(s804,s860,s776);
  nand x238(s806,s860,s780);
  nand x239(s855,s707,s721,s736);
  nand x240(s867,s707,s724,s736,s794);
  nand x241(s903,s3090,s3093);
  not x242(s3094,s3090);
  nand x243(s912,s3106,s3109);
  not x244(s3110,s3106);
  not x245(s915,s861);
  not x246(s927,s893);
  not x247(s941,s864);
  and x248(s977,s828,s974);
  and x249(s978,s150,s975);
  and x250(s984,s833,s981);
  and x251(s985,s159,s982);
  and x252(s991,s77,s988);
  and x253(s992,s50,s989);
  and x254(s998,s839,s995);
  and x255(s999,s828,s996);
  and x256(s1005,s845,s1002);
  and x257(s1006,s833,s1003);
  and x258(s1012,s107,s1009);
  and x259(s1013,s77,s1010);
  and x260(s1019,s116,s1016);
  and x261(s1020,s839,s1017);
  and x262(s1026,s283,s1023);
  and x263(s1027,s845,s1024);
  and x264(s1060,s200,s1054);
  and x265(s1063,s1048,s1054);
  and x266(s1066,s1049,s1057);
  and x267(s1069,s1050,s1057);
  nand x268(s1527,s784,s794);
  nand x269(s1530,s776,s794);
  nand x270(s1542,s707,s721,s1541);
  nand x271(s1563,s724,s732,s784);
  nand x272(s1572,s724,s784);
  not x273(s1581,s1512);
  not x274(s1585,s1512);
  not x275(s1589,s1512);
  not x276(s1593,s1512);
  not x277(s1597,s1512);
  not x278(s1601,s1512);
  not x279(s1605,s1512);
  not x280(s1716,s1681);
  and x281(s1718,s1681,s1699);
  not x282(s1723,s1681);
  and x283(s1725,s1681,s1699);
  not x284(s1730,s1681);
  and x285(s1732,s1681,s1699);
  not x286(s1737,s1681);
  and x287(s1739,s1681,s1699);
  not x288(s1744,s1681);
  and x289(s1746,s1681,s1699);
  not x290(s1751,s1681);
  and x291(s1753,s1681,s1699);
  not x292(s1758,s1681);
  and x293(s1760,s1681,s1699);
  not x294(s1765,s1681);
  and x295(s1767,s1681,s1699);
  and x296(s1852,s1834,s1773);
  nor x297(s1856,s50,s1773);
  not x298(s1870,s807);
  and x299(s1902,s1834,s1773);
  nor x300(s1906,s58,s1773);
  not x301(s1920,s807);
  and x302(s1953,s1834,s1773);
  nor x303(s1957,s68,s1773);
  not x304(s1971,s807);
  and x305(s2003,s1834,s1773);
  nor x306(s2007,s77,s1773);
  not x307(s2021,s807);
  and x308(s2058,s1834,s1773);
  nor x309(s2062,s87,s1773);
  not x310(s2076,s823);
  and x311(s2110,s1834,s1773);
  nor x312(s2114,s97,s1773);
  not x313(s2128,s816);
  and x314(s2163,s1834,s1773);
  nor x315(s2167,s107,s1773);
  not x316(s2181,s816);
  and x317(s2215,s1834,s1773);
  nor x318(s2219,s116,s1773);
  not x319(s2233,s816);
  and x320(s2285,s2278,s213);
  nand x321(s2288,s2278,s213);
  and x322(s2289,s2278,s213,s343);
  nand x323(s2293,s2278,s213,s343);
  and x324(s2298,s2278,s213,s343);
  nand x325(s2302,s2278,s213,s343);
  buf x326(s2877,s2874);
  nand x327(s2983,s2955,s2956);
  nand x328(s2986,s2965,s2966);
  not x329(s3014,s3010);
  nand x330(s3015,s3010,s3013);
  not x331(s3023,s3017);
  not x332(s3024,s3020);
  not x333(s3033,s3027);
  not x334(s3034,s3030);
  not x335(s3043,s3037);
  not x336(s3044,s3040);
  not x337(s355,s354);
  nand x338(s643,s3079,s3086);
  nand x339(s647,s3095,s3102);
  and x340(s680,s650,s675);
  nand x341(s904,s3087,s3094);
  nand x342(s913,s3103,s3110);
  and x343(s920,s588,s915);
  or x344(s979,s976,s977,s978);
  or x345(s993,s990,s991,s992);
  or x346(s1000,s997,s998,s999);
  or x347(s1007,s1004,s1005,s1006);
  or x348(s1021,s1018,s1019,s1020);
  or x349(s1028,s1025,s1026,s1027);
  and x350(s1719,s77,s1716);
  and x351(s1721,s223,s1718);
  and x352(s1726,s87,s1723);
  and x353(s1728,s226,s1725);
  and x354(s1733,s97,s1730);
  and x355(s1735,s232,s1732);
  and x356(s1740,s107,s1737);
  and x357(s1742,s238,s1739);
  and x358(s1747,s116,s1744);
  and x359(s1749,s244,s1746);
  and x360(s1754,s283,s1751);
  and x361(s1756,s250,s1753);
  and x362(s1761,s294,s1758);
  and x363(s1763,s257,s1760);
  and x364(s1768,s303,s1765);
  and x365(s1770,s264,s1767);
  buf x366(s1794,s1791);
  not x367(s1799,s1791);
  buf x368(s1812,s1809);
  not x369(s1817,s1809);
  and x370(s1859,s50,s1829,s1852);
  and x371(s1909,s58,s1829,s1902);
  and x372(s1960,s68,s1829,s1953);
  and x373(s2010,s77,s1829,s2003);
  and x374(s2065,s87,s2052,s2058);
  and x375(s2117,s97,s2052,s2110);
  and x376(s2170,s107,s2052,s2163);
  and x377(s2222,s116,s2052,s2215);
  not x378(s2678,s956);
  not x379(s2697,s956);
  not x380(s2716,s956);
  not x381(s2733,s956);
  not x382(s2751,s956);
  not x383(s2768,s956);
  not x384(s2785,s956);
  not x385(s2802,s956);
  nand x386(s3016,s3007,s3014);
  nand x387(s3025,s3020,s3023);
  nand x388(s3026,s3017,s3024);
  nand x389(s3035,s3030,s3033);
  nand x390(s3036,s3027,s3034);
  nand x391(s3045,s3040,s3043);
  nand x392(s3046,s3037,s3044);
  not x393(s2989,s2983);
  not x394(s2990,s2986);
  not x395(s610,s804);
  and x396(s613,s804,s806);
  not x397(s616,s806);
  nand x398(s640,s642,s643);
  nand x399(s648,s646,s647);
  and x400(s655,s630,s635,s442,s58);
  not x401(s665,s804);
  and x402(s668,s804,s806);
  not x403(s671,s806);
  not x404(s683,s804);
  not x405(s685,s806);
  and x406(s688,s804,s806);
  not x407(s694,s804);
  not x408(s696,s806);
  and x409(s699,s804,s806);
  buf x410(s870,s867);
  buf x411(s887,s867);
  nand x412(s901,s903,s904);
  nand x413(s910,s912,s913);
  not x414(s914,s855);
  and x415(s916,s855,s861);
  not x416(s942,s855);
  and x417(s943,s864,s855);
  nand x418(s1072,s1043,s1069);
  nand x419(s1084,s1043,s1066);
  nand x420(s1096,s1038,s1069);
  nand x421(s1108,s1038,s1066);
  nand x422(s1120,s1043,s1063);
  nand x423(s1132,s1043,s1060);
  nand x424(s1144,s1038,s1063);
  nand x425(s1156,s1038,s1060);
  not x426(s1533,s1527);
  not x427(s1534,s1530);
  and x428(s1535,s1527,s1530);
  buf x429(s1545,s1542);
  buf x430(s1554,s1542);
  not x431(s1610,s1572);
  not x432(s1619,s1572);
  not x433(s1628,s1572);
  not x434(s1637,s1572);
  not x435(s1646,s1563);
  not x436(s1655,s1563);
  not x437(s1664,s1563);
  not x438(s1673,s1563);
  or x439(s1722,s1719,s1720,s1721);
  or x440(s1729,s1726,s1727,s1728);
  or x441(s1736,s1733,s1734,s1735);
  or x442(s1743,s1740,s1741,s1742);
  or x443(s1750,s1747,s1748,s1749);
  or x444(s1757,s1754,s1755,s1756);
  or x445(s1764,s1761,s1762,s1763);
  or x446(s1771,s1768,s1769,s1770);
  and x447(s1853,s979,s1851);
  and x448(s1954,s993,s1952);
  and x449(s2004,s1000,s2002);
  and x450(s2059,s1007,s2057);
  and x451(s2164,s1021,s2162);
  and x452(s2216,s1028,s2214);
  buf x453(s2485,s2293);
  and x454(s2900,s2877,s2897);
  nand x455(s2903,s2877,s2897);
  buf x456(s2967,s557);
  buf x457(s2970,s562);
  buf x458(s2975,s557);
  buf x459(s2978,s562);
  nand x460(s3047,s3015,s3016);
  nand x461(s3050,s3025,s3026);
  nand x462(s3055,s3035,s3036);
  nand x463(s3058,s3045,s3046);
  nand x464(s574,s2986,s2989);
  nand x465(s575,s2983,s2990);
  and x466(s617,s501,s613);
  and x467(s641,s640,s476,s639);
  and x468(s649,s530,s648);
  and x469(s662,s655,s657);
  and x470(s672,s513,s668);
  and x471(s690,s654,s685);
  and x472(s691,s540,s688);
  and x473(s701,s634,s696);
  and x474(s702,s526,s699);
  not x475(s902,s901);
  not x476(s911,s910);
  and x477(s917,s650,s914);
  and x478(s923,s586,s916);
  and x479(s1538,s442,s1535);
  and x480(s1871,s1817,s226,s1870);
  and x481(s1872,s1817,s274,s807);
  and x482(s1873,s1812,s1722);
  and x483(s1921,s1817,s232,s1920);
  and x484(s1922,s1817,s274,s807);
  and x485(s1923,s1812,s1729);
  and x486(s1972,s1817,s238,s1971);
  and x487(s1973,s1817,s274,s807);
  and x488(s1974,s1812,s1736);
  and x489(s2022,s1817,s244,s2021);
  and x490(s2023,s1817,s274,s807);
  and x491(s2024,s1812,s1743);
  and x492(s2077,s1799,s250,s2076);
  and x493(s2078,s1799,s274,s823);
  and x494(s2079,s1794,s1750);
  and x495(s2129,s1799,s257,s2128);
  and x496(s2130,s1799,s274,s816);
  and x497(s2131,s1794,s1757);
  and x498(s2182,s1799,s264,s2181);
  and x499(s2183,s1799,s274,s816);
  and x500(s2184,s1794,s1764);
  and x501(s2234,s1799,s270,s2233);
  and x502(s2235,s1799,s274,s816);
  and x503(s2236,s1794,s1771);
  not x504(s2973,s2967);
  not x505(s2974,s2970);
  not x506(s2981,s2975);
  not x507(s2982,s2978);
  nand x508(s576,s574,s575);
  not x509(s3053,s3047);
  not x510(s3054,s3050);
  not x511(s3061,s3055);
  not x512(s3062,s3058);
  or x513(s645,s641,s644);
  not x514(s926,s887);
  and x515(s928,s887,s893);
  and x516(s947,s649,s942);
  and x517(s983,s902,s980);
  and x518(s1011,s911,s1008);
  buf x519(s1075,s1072);
  buf x520(s1087,s1084);
  buf x521(s1099,s1096);
  buf x522(s1111,s1108);
  buf x523(s1123,s1120);
  buf x524(s1135,s1132);
  buf x525(s1147,s1144);
  buf x526(s1159,s1156);
  buf x527(s1168,s1072);
  buf x528(s1177,s1084);
  buf x529(s1186,s1096);
  buf x530(s1195,s1108);
  buf x531(s1204,s1120);
  buf x532(s1213,s1132);
  buf x533(s1222,s1144);
  buf x534(s1231,s1156);
  not x535(s1609,s1545);
  and x536(s1611,s1545,s1572);
  not x537(s1618,s1545);
  and x538(s1620,s1545,s1572);
  not x539(s1627,s1545);
  and x540(s1629,s1545,s1572);
  not x541(s1636,s1545);
  and x542(s1638,s1545,s1572);
  not x543(s1645,s1554);
  and x544(s1647,s1554,s1563);
  not x545(s1654,s1554);
  and x546(s1656,s1554,s1563);
  not x547(s1663,s1554);
  and x548(s1665,s1554,s1563);
  not x549(s1672,s1554);
  and x550(s1674,s1554,s1563);
  or x551(s1862,s1853,s1856,s1859);
  nor x552(s1866,s1853,s1856,s1859);
  or x553(s1874,s1871,s1872,s1873);
  or x554(s1924,s1921,s1922,s1923);
  or x555(s1963,s1954,s1957,s1960);
  nor x556(s1967,s1954,s1957,s1960);
  or x557(s1975,s1972,s1973,s1974);
  or x558(s2013,s2004,s2007,s2010);
  nor x559(s2017,s2004,s2007,s2010);
  or x560(s2025,s2022,s2023,s2024);
  or x561(s2068,s2059,s2062,s2065);
  nor x562(s2072,s2059,s2062,s2065);
  or x563(s2080,s2077,s2078,s2079);
  or x564(s2132,s2129,s2130,s2131);
  or x565(s2173,s2164,s2167,s2170);
  nor x566(s2177,s2164,s2167,s2170);
  or x567(s2185,s2182,s2183,s2184);
  or x568(s2225,s2216,s2219,s2222);
  nor x569(s2229,s2216,s2219,s2222);
  or x570(s2237,s2234,s2235,s2236);
  not x571(s2488,s2485);
  not x572(s2679,s870);
  and x573(s2680,s956,s870);
  not x574(s2698,s870);
  and x575(s2699,s956,s870);
  not x576(s2717,s870);
  and x577(s2718,s956,s870);
  not x578(s2734,s870);
  and x579(s2735,s956,s870);
  not x580(s2752,s870);
  and x581(s2753,s956,s870);
  not x582(s2769,s870);
  and x583(s2770,s956,s870);
  not x584(s2786,s870);
  and x585(s2787,s956,s870);
  not x586(s2803,s870);
  and x587(s2804,s956,s870);
  or x588(s359,s917,s920,s923);
  nor x589(s1029,s917,s920,s923);
  nand x590(s565,s2970,s2973);
  nand x591(s566,s2967,s2974);
  nand x592(s569,s2978,s2981);
  nand x593(s570,s2975,s2982);
  nand x594(s589,s3050,s3053);
  nand x595(s590,s3047,s3054);
  nand x596(s595,s3058,s3061);
  nand x597(s596,s3055,s3062);
  and x598(s929,s650,s926);
  and x599(s938,s630,s928);
  and x600(s944,s645,s941);
  or x601(s986,s983,s984,s985);
  or x602(s1014,s1011,s1012,s1013);
  and x603(s1616,s442,s1611);
  and x604(s1625,s456,s1620);
  and x605(s1634,s463,s1629);
  and x606(s1643,s479,s1638);
  not x607(s360,s1029);
  nand x608(s567,s565,s566);
  nand x609(s571,s569,s570);
  buf x610(s579,s576);
  nand x611(s591,s589,s590);
  nand x612(s597,s595,s596);
  and x613(s614,s576,s610);
  not x614(s1240,s1075);
  not x615(s1241,s1087);
  not x616(s1242,s1099);
  not x617(s1243,s1111);
  not x618(s1244,s1123);
  not x619(s1245,s1135);
  not x620(s1246,s1147);
  not x621(s1247,s1159);
  not x622(s1257,s1075);
  not x623(s1258,s1087);
  not x624(s1259,s1099);
  not x625(s1260,s1111);
  not x626(s1261,s1123);
  not x627(s1262,s1135);
  not x628(s1263,s1147);
  not x629(s1264,s1159);
  not x630(s1274,s1075);
  not x631(s1275,s1087);
  not x632(s1276,s1099);
  not x633(s1277,s1111);
  not x634(s1278,s1123);
  not x635(s1279,s1135);
  not x636(s1280,s1147);
  not x637(s1281,s1159);
  not x638(s1291,s1075);
  not x639(s1292,s1087);
  not x640(s1293,s1099);
  not x641(s1294,s1111);
  not x642(s1295,s1123);
  not x643(s1296,s1135);
  not x644(s1297,s1147);
  not x645(s1298,s1159);
  not x646(s1308,s1075);
  not x647(s1309,s1087);
  not x648(s1310,s1099);
  not x649(s1311,s1111);
  not x650(s1312,s1123);
  not x651(s1313,s1135);
  not x652(s1314,s1147);
  not x653(s1315,s1159);
  not x654(s1325,s1075);
  not x655(s1326,s1087);
  not x656(s1327,s1099);
  not x657(s1328,s1111);
  not x658(s1329,s1123);
  not x659(s1330,s1135);
  not x660(s1331,s1147);
  not x661(s1332,s1159);
  not x662(s1342,s1075);
  not x663(s1343,s1087);
  not x664(s1344,s1099);
  not x665(s1345,s1111);
  not x666(s1346,s1123);
  not x667(s1347,s1135);
  not x668(s1348,s1147);
  not x669(s1349,s1159);
  not x670(s1359,s1075);
  not x671(s1360,s1087);
  not x672(s1361,s1099);
  not x673(s1362,s1111);
  not x674(s1363,s1123);
  not x675(s1364,s1135);
  not x676(s1365,s1147);
  not x677(s1366,s1159);
  not x678(s1376,s1168);
  not x679(s1377,s1177);
  not x680(s1378,s1186);
  not x681(s1379,s1195);
  not x682(s1380,s1204);
  not x683(s1381,s1213);
  not x684(s1382,s1222);
  not x685(s1383,s1231);
  not x686(s1393,s1168);
  not x687(s1394,s1177);
  not x688(s1395,s1186);
  not x689(s1396,s1195);
  not x690(s1397,s1204);
  not x691(s1398,s1213);
  not x692(s1399,s1222);
  not x693(s1400,s1231);
  not x694(s1410,s1168);
  not x695(s1411,s1177);
  not x696(s1412,s1186);
  not x697(s1413,s1195);
  not x698(s1414,s1204);
  not x699(s1415,s1213);
  not x700(s1416,s1222);
  not x701(s1417,s1231);
  not x702(s1427,s1168);
  not x703(s1428,s1177);
  not x704(s1429,s1186);
  not x705(s1430,s1195);
  not x706(s1431,s1204);
  not x707(s1432,s1213);
  not x708(s1433,s1222);
  not x709(s1434,s1231);
  not x710(s1444,s1168);
  not x711(s1445,s1177);
  not x712(s1446,s1186);
  not x713(s1447,s1195);
  not x714(s1448,s1204);
  not x715(s1449,s1213);
  not x716(s1450,s1222);
  not x717(s1451,s1231);
  not x718(s1461,s1168);
  not x719(s1462,s1177);
  not x720(s1463,s1186);
  not x721(s1464,s1195);
  not x722(s1465,s1204);
  not x723(s1466,s1213);
  not x724(s1467,s1222);
  not x725(s1468,s1231);
  not x726(s1478,s1168);
  not x727(s1479,s1177);
  not x728(s1480,s1186);
  not x729(s1481,s1195);
  not x730(s1482,s1204);
  not x731(s1483,s1213);
  not x732(s1484,s1222);
  not x733(s1485,s1231);
  not x734(s1495,s1168);
  not x735(s1496,s1177);
  not x736(s1497,s1186);
  not x737(s1498,s1195);
  not x738(s1499,s1204);
  not x739(s1500,s1213);
  not x740(s1501,s1222);
  not x741(s1502,s1231);
  buf x742(s1877,s1874);
  not x743(s1880,s1874);
  not x744(s1891,s1866);
  and x745(s1903,s986,s1901);
  buf x746(s1927,s1924);
  not x747(s1930,s1924);
  buf x748(s1978,s1975);
  not x749(s1981,s1975);
  not x750(s1992,s1967);
  buf x751(s2028,s2025);
  not x752(s2031,s2025);
  not x753(s2042,s2017);
  buf x754(s2085,s2080);
  not x755(s2088,s2080);
  not x756(s2099,s2072);
  and x757(s2111,s1014,s2109);
  buf x758(s2137,s2132);
  not x759(s2140,s2132);
  buf x760(s2190,s2185);
  not x761(s2193,s2185);
  not x762(s2204,s2177);
  buf x763(s2242,s2237);
  not x764(s2245,s2237);
  not x765(s2256,s2229);
  and x766(s2320,s2285,s1862);
  and x767(s2341,s2289,s1963);
  and x768(s2354,s2289,s2013);
  and x769(s2367,s2289,s2068);
  and x770(s2383,s2298,s2173);
  and x771(s2391,s2298,s2225);
  not x772(s2474,s2080);
  not x773(s2475,s2132);
  not x774(s2476,s2185);
  not x775(s2477,s2237);
  and x776(s2482,s2080,s2132,s2185,s2237,s2481);
  nand x777(s361,s359,s360);
  not x778(s568,s567);
  or x779(s618,s614,s616,s617);
  and x780(s1248,s124,s1240);
  and x781(s1249,s159,s1241);
  and x782(s1250,s150,s1242);
  and x783(s1251,s143,s1243);
  and x784(s1252,s137,s1244);
  and x785(s1253,s132,s1245);
  and x786(s1254,s128,s1246);
  and x787(s1255,s125,s1247);
  and x788(s1265,s125,s1257);
  and x789(s1266,s432,s1258);
  and x790(s1267,s159,s1259);
  and x791(s1268,s150,s1260);
  and x792(s1269,s143,s1261);
  and x793(s1270,s137,s1262);
  and x794(s1271,s132,s1263);
  and x795(s1272,s128,s1264);
  and x796(s1282,s128,s1274);
  and x797(s1283,s447,s1275);
  and x798(s1284,s432,s1276);
  and x799(s1285,s159,s1277);
  and x800(s1286,s150,s1278);
  and x801(s1287,s143,s1279);
  and x802(s1288,s137,s1280);
  and x803(s1289,s132,s1281);
  and x804(s1299,s132,s1291);
  and x805(s1300,s467,s1292);
  and x806(s1301,s447,s1293);
  and x807(s1302,s432,s1294);
  and x808(s1303,s159,s1295);
  and x809(s1304,s150,s1296);
  and x810(s1305,s143,s1297);
  and x811(s1306,s137,s1298);
  and x812(s1316,s137,s1308);
  and x813(s1317,s483,s1309);
  and x814(s1318,s467,s1310);
  and x815(s1319,s447,s1311);
  and x816(s1320,s432,s1312);
  and x817(s1321,s159,s1313);
  and x818(s1322,s150,s1314);
  and x819(s1323,s143,s1315);
  and x820(s1333,s143,s1325);
  and x821(s1334,s492,s1326);
  and x822(s1335,s483,s1327);
  and x823(s1336,s467,s1328);
  and x824(s1337,s447,s1329);
  and x825(s1338,s432,s1330);
  and x826(s1339,s159,s1331);
  and x827(s1340,s150,s1332);
  and x828(s1350,s150,s1342);
  and x829(s1351,s504,s1343);
  and x830(s1352,s492,s1344);
  and x831(s1353,s483,s1345);
  and x832(s1354,s467,s1346);
  and x833(s1355,s447,s1347);
  and x834(s1356,s432,s1348);
  and x835(s1357,s159,s1349);
  and x836(s1367,s159,s1359);
  and x837(s1368,s517,s1360);
  and x838(s1369,s504,s1361);
  and x839(s1370,s492,s1362);
  and x840(s1371,s483,s1363);
  and x841(s1372,s467,s1364);
  and x842(s1373,s447,s1365);
  and x843(s1374,s432,s1366);
  and x844(s1384,s283,s1376);
  and x845(s1385,s447,s1377);
  and x846(s1386,s467,s1378);
  and x847(s1387,s483,s1379);
  and x848(s1388,s492,s1380);
  and x849(s1389,s504,s1381);
  and x850(s1390,s517,s1382);
  and x851(s1391,s530,s1383);
  and x852(s1401,s294,s1393);
  and x853(s1402,s467,s1394);
  and x854(s1403,s483,s1395);
  and x855(s1404,s492,s1396);
  and x856(s1405,s504,s1397);
  and x857(s1406,s517,s1398);
  and x858(s1407,s530,s1399);
  and x859(s1408,s283,s1400);
  and x860(s1418,s303,s1410);
  and x861(s1419,s483,s1411);
  and x862(s1420,s492,s1412);
  and x863(s1421,s504,s1413);
  and x864(s1422,s517,s1414);
  and x865(s1423,s530,s1415);
  and x866(s1424,s283,s1416);
  and x867(s1425,s294,s1417);
  and x868(s1435,s311,s1427);
  and x869(s1436,s492,s1428);
  and x870(s1437,s504,s1429);
  and x871(s1438,s517,s1430);
  and x872(s1439,s530,s1431);
  and x873(s1440,s283,s1432);
  and x874(s1441,s294,s1433);
  and x875(s1442,s303,s1434);
  and x876(s1452,s317,s1444);
  and x877(s1453,s504,s1445);
  and x878(s1454,s517,s1446);
  and x879(s1455,s530,s1447);
  and x880(s1456,s283,s1448);
  and x881(s1457,s294,s1449);
  and x882(s1458,s303,s1450);
  and x883(s1459,s311,s1451);
  and x884(s1469,s322,s1461);
  and x885(s1470,s517,s1462);
  and x886(s1471,s530,s1463);
  and x887(s1472,s283,s1464);
  and x888(s1473,s294,s1465);
  and x889(s1474,s303,s1466);
  and x890(s1475,s311,s1467);
  and x891(s1476,s317,s1468);
  and x892(s1486,s326,s1478);
  and x893(s1487,s530,s1479);
  and x894(s1488,s283,s1480);
  and x895(s1489,s294,s1481);
  and x896(s1490,s303,s1482);
  and x897(s1491,s311,s1483);
  and x898(s1492,s317,s1484);
  and x899(s1493,s322,s1485);
  and x900(s1503,s329,s1495);
  and x901(s1504,s283,s1496);
  and x902(s1505,s294,s1497);
  and x903(s1506,s303,s1498);
  and x904(s1507,s311,s1499);
  and x905(s1508,s317,s1500);
  and x906(s1509,s322,s1501);
  and x907(s1510,s326,s1502);
  and x908(s2483,s2474,s2475,s2476,s2477,s2478);
  buf x909(s600,s597);
  and x910(s661,s568,s660);
  and x911(s669,s597,s665);
  and x912(s679,s591,s678);
  nor x913(s1256,s1248,s1249,s1250,s1251,s1252,s1253,s1254,s1255);
  nor x914(s1273,s1265,s1266,s1267,s1268,s1269,s1270,s1271,s1272);
  nor x915(s1290,s1282,s1283,s1284,s1285,s1286,s1287,s1288,s1289);
  nor x916(s1307,s1299,s1300,s1301,s1302,s1303,s1304,s1305,s1306);
  nor x917(s1324,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323);
  nor x918(s1341,s1333,s1334,s1335,s1336,s1337,s1338,s1339,s1340);
  nor x919(s1358,s1350,s1351,s1352,s1353,s1354,s1355,s1356,s1357);
  nor x920(s1375,s1367,s1368,s1369,s1370,s1371,s1372,s1373,s1374);
  nor x921(s1392,s1384,s1385,s1386,s1387,s1388,s1389,s1390,s1391);
  nor x922(s1409,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408);
  nor x923(s1426,s1418,s1419,s1420,s1421,s1422,s1423,s1424,s1425);
  nor x924(s1443,s1435,s1436,s1437,s1438,s1439,s1440,s1441,s1442);
  nor x925(s1460,s1452,s1453,s1454,s1455,s1456,s1457,s1458,s1459);
  nor x926(s1477,s1469,s1470,s1471,s1472,s1473,s1474,s1475,s1476);
  nor x927(s1494,s1486,s1487,s1488,s1489,s1490,s1491,s1492,s1493);
  nor x928(s1511,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510);
  and x929(s1652,s618,s1647);
  and x930(s1883,s169,s1862,s1877);
  and x931(s1886,s179,s1862,s1880);
  and x932(s1889,s190,s1866,s1880);
  and x933(s1890,s200,s1866,s1877);
  or x934(s1912,s1903,s1906,s1909);
  nor x935(s1916,s1903,s1906,s1909);
  and x936(s1984,s169,s1963,s1978);
  and x937(s1987,s179,s1963,s1981);
  and x938(s1990,s190,s1967,s1981);
  and x939(s1991,s200,s1967,s1978);
  and x940(s2034,s169,s2013,s2028);
  and x941(s2037,s179,s2013,s2031);
  and x942(s2040,s190,s2017,s2031);
  and x943(s2041,s200,s2017,s2028);
  and x944(s2091,s169,s2068,s2085);
  and x945(s2094,s179,s2068,s2088);
  and x946(s2097,s190,s2072,s2088);
  and x947(s2098,s200,s2072,s2085);
  or x948(s2120,s2111,s2114,s2117);
  nor x949(s2124,s2111,s2114,s2117);
  and x950(s2196,s169,s2173,s2190);
  and x951(s2199,s179,s2173,s2193);
  and x952(s2202,s190,s2177,s2193);
  and x953(s2203,s200,s2177,s2190);
  and x954(s2248,s169,s2225,s2242);
  and x955(s2251,s179,s2225,s2245);
  and x956(s2254,s190,s2229,s2245);
  and x957(s2255,s200,s2229,s2242);
  or x958(s2484,s2482,s2483);
  buf x959(s2991,s571);
  buf x960(s2994,s579);
  buf x961(s2999,s571);
  buf x962(s3002,s579);
  buf x963(s3063,s591);
  buf x964(s3071,s591);
  buf x965(s3124,s2320);
  buf x966(s3134,s2320);
  buf x967(s3158,s2341);
  buf x968(s3166,s2341);
  buf x969(s3174,s2354);
  buf x970(s3182,s2354);
  buf x971(s3190,s2367);
  buf x972(s3200,s2367);
  buf x973(s3224,s2383);
  buf x974(s3232,s2383);
  buf x975(s3240,s2391);
  buf x976(s3248,s2391);
  nor x977(s663,s661,s662);
  or x978(s673,s669,s671,s672);
  nor x979(s681,s679,s680);
  and x980(s1536,s1256,s1533);
  and x981(s1537,s1392,s1534);
  and x982(s1582,s1273,s1581);
  and x983(s1583,s1409,s1512);
  and x984(s1586,s1290,s1585);
  and x985(s1587,s1426,s1512);
  and x986(s1590,s1307,s1589);
  and x987(s1591,s1443,s1512);
  and x988(s1594,s1324,s1593);
  and x989(s1595,s1460,s1512);
  and x990(s1598,s1341,s1597);
  and x991(s1599,s1477,s1512);
  and x992(s1602,s1358,s1601);
  and x993(s1603,s1494,s1512);
  and x994(s1606,s1375,s1605);
  and x995(s1607,s1511,s1512);
  or x996(s1894,s1889,s1890,s1891);
  or x997(s1997,s1990,s1991,s1992);
  or x998(s2047,s2040,s2041,s2042);
  or x999(s2102,s2097,s2098,s2099);
  or x1000(s2209,s2202,s2203,s2204);
  or x1001(s2261,s2254,s2255,s2256);
  and x1002(s2489,s2484,s2488);
  not x1003(s3005,s2999);
  not x1004(s3006,s3002);
  not x1005(s3077,s3071);
  not x1006(s3069,s3063);
  not x1007(s2997,s2991);
  not x1008(s2998,s2994);
  and x1009(s689,s681,s683);
  and x1010(s700,s663,s694);
  or x1011(s1539,s1536,s1537,s1538);
  or x1012(s1584,s1582,s1583);
  or x1013(s1588,s1586,s1587);
  or x1014(s1592,s1590,s1591);
  or x1015(s1596,s1594,s1595);
  or x1016(s1600,s1598,s1599);
  or x1017(s1604,s1602,s1603);
  or x1018(s1608,s1606,s1607);
  and x1019(s1661,s673,s1656);
  or x1020(s1892,s1883,s1886);
  nor x1021(s1893,s1883,s1886);
  and x1022(s1933,s169,s1912,s1927);
  and x1023(s1936,s179,s1912,s1930);
  and x1024(s1939,s190,s1916,s1930);
  and x1025(s1940,s200,s1916,s1927);
  not x1026(s1941,s1916);
  or x1027(s1993,s1984,s1987);
  nor x1028(s1996,s1984,s1987);
  or x1029(s2043,s2034,s2037);
  nor x1030(s2046,s2034,s2037);
  or x1031(s2100,s2091,s2094);
  nor x1032(s2101,s2091,s2094);
  and x1033(s2143,s169,s2120,s2137);
  and x1034(s2146,s179,s2120,s2140);
  and x1035(s2149,s190,s2124,s2140);
  and x1036(s2150,s200,s2124,s2137);
  not x1037(s2151,s2124);
  or x1038(s2205,s2196,s2199);
  nor x1039(s2208,s2196,s2199);
  or x1040(s2257,s2248,s2251);
  nor x1041(s2260,s2248,s2251);
  not x1042(s3138,s3134);
  and x1043(s2328,s2285,s1912);
  not x1044(s3162,s3158);
  not x1045(s3170,s3166);
  not x1046(s3178,s3174);
  not x1047(s3186,s3182);
  not x1048(s3204,s3200);
  and x1049(s2375,s2298,s2120);
  not x1050(s3236,s3232);
  not x1051(s3244,s3240);
  not x1052(s3252,s3248);
  not x1053(s3228,s3224);
  buf x1054(s3066,s600);
  buf x1055(s3074,s600);
  not x1056(s3128,s3124);
  not x1057(s3194,s3190);
  nand x1058(s619,s2994,s2997);
  nand x1059(s620,s2991,s2998);
  nand x1060(s582,s3002,s3005);
  nand x1061(s583,s2999,s3006);
  or x1062(s692,s689,s690,s691);
  or x1063(s703,s700,s701,s702);
  and x1064(s1612,s1539,s1609);
  and x1065(s1621,s1584,s1618);
  and x1066(s1630,s1588,s1627);
  and x1067(s1639,s1592,s1636);
  and x1068(s1648,s1596,s1645);
  and x1069(s1657,s1600,s1654);
  and x1070(s1666,s1604,s1663);
  and x1071(s1675,s1608,s1672);
  and x1072(s1895,s1893,s1894);
  or x1073(s1946,s1939,s1940,s1941);
  and x1074(s1998,s1996,s1997);
  and x1075(s2048,s2046,s2047);
  and x1076(s2103,s2101,s2102);
  or x1077(s2156,s2149,s2150,s2151);
  and x1078(s2210,s2208,s2209);
  and x1079(s2262,s2260,s2261);
  not x1080(s2271,s1892);
  not x1081(s2311,s2100);
  nand x1082(s356,s619,s620);
  nand x1083(s357,s582,s583);
  nand x1084(s603,s3074,s3077);
  not x1085(s3078,s3074);
  nand x1086(s606,s3066,s3069);
  not x1087(s3070,s3066);
  and x1088(s1670,s703,s1665);
  and x1089(s1679,s692,s1674);
  or x1090(s1942,s1933,s1936);
  nor x1091(s1945,s1933,s1936);
  or x1092(s2152,s2143,s2146);
  nor x1093(s2155,s2143,s2146);
  and x1094(s2445,s1993,s2293);
  and x1095(s2448,s2043,s2293);
  and x1096(s2455,s2205,s2302);
  and x1097(s2458,s2257,s2302);
  buf x1098(s3142,s2328);
  buf x1099(s3150,s2328);
  buf x1100(s3208,s2375);
  buf x1101(s3216,s2375);
  nand x1102(s358,s356,s357);
  nand x1103(s604,s3071,s3078);
  nand x1104(s607,s3063,s3070);
  and x1105(s1947,s1945,s1946);
  and x1106(s2157,s2155,s2156);
  buf x1107(s2317,s1895);
  buf x1108(s2338,s1998);
  buf x1109(s2351,s2048);
  buf x1110(s2364,s2103);
  buf x1111(s2380,s2210);
  buf x1112(s2388,s2262);
  nand x1113(s605,s603,s604);
  nand x1114(s608,s606,s607);
  nand x1115(s2272,s1895,s1942);
  nand x1116(s2312,s2103,s2152);
  not x1117(s3146,s3142);
  not x1118(s3154,s3150);
  not x1119(s3220,s3216);
  not x1120(s3212,s3208);
  and x1121(s2444,s1942,s2288);
  buf x1122(s2451,s2448);
  and x1123(s2454,s2152,s2293);
  buf x1124(s2461,s2458);
  not x1125(s2530,s2445);
  buf x1126(s3323,s2458);
  not x1127(s349,s605);
  not x1128(s350,s608);
  and x1129(s2265,s1895,s1947,s1998,s2048);
  nand x1130(s2273,s1895,s1947,s1993);
  nand x1131(s2274,s2043,s1947,s1998,s1895);
  and x1132(s2309,s2103,s2157,s2210,s2262);
  nand x1133(s2313,s2103,s2157,s2205);
  nand x1134(s2314,s2257,s2157,s2210,s2103);
  buf x1135(s2325,s1947);
  buf x1136(s2372,s2157);
  not x1137(s2523,s2444);
  not x1138(s2533,s2454);
  buf x1139(s3121,s2317);
  buf x1140(s3131,s2317);
  buf x1141(s3155,s2338);
  buf x1142(s3163,s2338);
  buf x1143(s3171,s2351);
  buf x1144(s3179,s2351);
  buf x1145(s3187,s2364);
  buf x1146(s3197,s2364);
  buf x1147(s3221,s2380);
  buf x1148(s3229,s2380);
  buf x1149(s3237,s2388);
  buf x1150(s3245,s2388);
  nand x1151(s351,s349,s350);
  nand x1152(s2275,s2271,s2272,s2273,s2274);
  nand x1153(s2315,s2311,s2312,s2313,s2314);
  not x1154(s3329,s3323);
  and x1155(s372,s2309,s2265);
  nand x1156(s2324,s3131,s3138);
  nand x1157(s2350,s3163,s3170);
  nand x1158(s2363,s3179,s3186);
  nand x1159(s2371,s3197,s3204);
  nand x1160(s2387,s3229,s3236);
  nand x1161(s2400,s3245,s3252);
  buf x1162(s2268,s2265);
  not x1163(s3137,s3131);
  not x1164(s3161,s3155);
  nand x1165(s2345,s3155,s3162);
  not x1166(s3169,s3163);
  not x1167(s3177,s3171);
  nand x1168(s2358,s3171,s3178);
  not x1169(s3185,s3179);
  not x1170(s3203,s3197);
  not x1171(s3235,s3229);
  not x1172(s3243,s3237);
  nand x1173(s2395,s3237,s3244);
  not x1174(s3251,s3245);
  not x1175(s3227,s3221);
  nand x1176(s2432,s3221,s3228);
  and x1177(s2490,s2309,s2485);
  not x1178(s3127,s3121);
  nand x1179(s3130,s3121,s3128);
  buf x1180(s3139,s2325);
  buf x1181(s3147,s2325);
  not x1182(s3193,s3187);
  nand x1183(s3196,s3187,s3194);
  buf x1184(s3205,s2372);
  buf x1185(s3213,s2372);
  nand x1186(s2307,s2265,s2315);
  not x1187(s2308,s2275);
  nand x1188(s2323,s3134,s3137);
  nand x1189(s2349,s3166,s3169);
  nand x1190(s2362,s3182,s3185);
  nand x1191(s2370,s3200,s3203);
  nand x1192(s2386,s3232,s3235);
  nand x1193(s2399,s3248,s3251);
  nand x1194(s2344,s3158,s3161);
  nand x1195(s2357,s3174,s3177);
  nand x1196(s2394,s3240,s3243);
  nand x1197(s2431,s3224,s3227);
  and x1198(s2464,s2315,s2302);
  or x1199(s2491,s2489,s2490);
  nand x1200(s3129,s3124,s3127);
  nand x1201(s3195,s3190,s3193);
  and x1202(s368,s2307,s2308);
  nand x1203(s1615,s2323,s2324);
  nand x1204(s2337,s3147,s3154);
  nand x1205(s1633,s2349,s2350);
  nand x1206(s1642,s2362,s2363);
  nand x1207(s1651,s2370,s2371);
  nand x1208(s2379,s3213,s3220);
  nand x1209(s1669,s2386,s2387);
  nand x1210(s1678,s2399,s2400);
  not x1211(s3145,s3139);
  nand x1212(s2332,s3139,s3146);
  not x1213(s3153,s3147);
  nand x1214(s2346,s2344,s2345);
  nand x1215(s2359,s2357,s2358);
  not x1216(s3219,s3213);
  nand x1217(s2396,s2394,s2395);
  not x1218(s3211,s3205);
  nand x1219(s2425,s3205,s3212);
  nand x1220(s2433,s2431,s2432);
  nand x1221(s3272,s3129,s3130);
  nand x1222(s3308,s3195,s3196);
  not x1223(s369,s368);
  not x1224(s1613,s1615);
  nand x1225(s2336,s3150,s3153);
  not x1226(s1631,s1633);
  not x1227(s1640,s1642);
  not x1228(s1649,s1651);
  nand x1229(s2378,s3216,s3219);
  not x1230(s1667,s1669);
  not x1231(s1676,s1678);
  nand x1232(s2331,s3142,s3145);
  nand x1233(s2424,s3208,s3211);
  buf x1234(s2467,s2464);
  buf x1235(s2495,s2491);
  buf x1236(s3295,s2464);
  and x1237(s3374,s330,s2491);
  and x1238(s1614,s1613,s1610);
  nand x1239(s1624,s2336,s2337);
  and x1240(s1632,s1631,s1628);
  and x1241(s1641,s1640,s1637);
  and x1242(s1650,s1649,s1646);
  nand x1243(s1660,s2378,s2379);
  and x1244(s1668,s1667,s1664);
  and x1245(s1677,s1676,s1673);
  nand x1246(s2333,s2331,s2332);
  buf x1247(s2406,s2346);
  buf x1248(s2409,s2346);
  buf x1249(s2415,s2359);
  buf x1250(s2419,s2359);
  nand x1251(s2426,s2424,s2425);
  buf x1252(s2439,s2396);
  and x1253(s2518,s2433,s2461);
  not x1254(s3276,s3272);
  not x1255(s3312,s3308);
  and x1256(s2612,s330,s2396);
  buf x1257(s3326,s2433);
  nor x1258(s1617,s1612,s1614,s1616);
  not x1259(s1622,s1624);
  nor x1260(s1635,s1630,s1632,s1634);
  nor x1261(s1644,s1639,s1641,s1643);
  nor x1262(s1653,s1648,s1650,s1652);
  not x1263(s1658,s1660);
  nor x1264(s1671,s1666,s1668,s1670);
  nor x1265(s1680,s1675,s1677,s1679);
  and x1266(s2500,s2467,s2268);
  and x1267(s2505,s2495,s2268);
  or x1268(s2519,s2455,s2518);
  not x1269(s3378,s3374);
  not x1270(s2642,s2467);
  buf x1271(s2645,s2467);
  not x1272(s3301,s3295);
  and x1273(s1623,s1622,s1619);
  and x1274(s1659,s1658,s1655);
  buf x1275(s2401,s2333);
  or x1276(s2501,s2275,s2500);
  and x1277(s2511,s2495,s2419,s2409);
  and x1278(s2512,s2495,s2415);
  and x1279(s2513,s2439,s2433,s2426);
  and x1280(s2514,s2439,s2433);
  and x1281(s2517,s2467,s2415);
  nand x1282(s2531,s2409,s2451);
  nand x1283(s2532,s2409,s2419,s2467);
  nand x1284(s2534,s2426,s2455);
  nand x1285(s2535,s2426,s2433,s2461);
  nand x1286(s2607,s3326,s3329);
  not x1287(s3330,s3326);
  and x1288(s2643,s330,s2491,s2642);
  and x1289(s2687,s1617,s2680);
  and x1290(s2725,s1635,s2718);
  and x1291(s2742,s1644,s2735);
  and x1292(s2760,s1653,s2753);
  and x1293(s2794,s1671,s2787);
  and x1294(s2811,s1680,s2804);
  buf x1295(s3280,s2333);
  buf x1296(s3290,s2409);
  buf x1297(s3298,s2415);
  buf x1298(s3316,s2426);
  buf x1299(s3406,s2612);
  buf x1300(s3414,s2612);
  and x1301(s3422,s2439,s2439);
  nor x1302(s1626,s1621,s1623,s1625);
  nor x1303(s1662,s1657,s1659,s1661);
  and x1304(s2567,s330,s2512);
  and x1305(s2589,s330,s2513);
  nand x1306(s2608,s3323,s3330);
  buf x1307(s2654,s2519);
  buf x1308(s3253,s2505);
  nand x1309(s3277,s2530,s2531,s2532);
  or x1310(s3287,s2448,s2517);
  nand x1311(s3305,s2533,s2534,s2535);
  buf x1312(s3313,s2519);
  and x1313(s3350,s330,s2511);
  or x1314(s932,s2643,s2645);
  and x1315(s2508,s2495,s2401,s2409,s2419);
  nand x1316(s2524,s2401,s2445);
  nand x1317(s2525,s2401,s2406,s2451);
  nand x1318(s2526,s2401,s2406,s2419,s2467);
  not x1319(s3294,s3290);
  nand x1320(s2609,s2607,s2608);
  not x1321(s3410,s3406);
  not x1322(s3418,s3414);
  nand x1323(s2624,s3422,s3425);
  not x1324(s3426,s3422);
  buf x1325(s2629,s2501);
  nor x1326(s2647,s2643,s2645);
  and x1327(s2706,s1626,s2699);
  and x1328(s2777,s1662,s2770);
  buf x1329(s3264,s2501);
  not x1330(s3284,s3280);
  not x1331(s3302,s3298);
  nand x1332(s3303,s3298,s3301);
  not x1333(s3320,s3316);
  and x1334(s3398,s330,s2514);
  not x1335(s2657,s2654);
  and x1336(s398,s2519,s2654);
  and x1337(s933,s932,s927);
  nand x1338(s2527,s2523,s2524,s2525,s2526);
  not x1339(s3259,s3253);
  not x1340(s3354,s3350);
  not x1341(s3293,s3287);
  nand x1342(s2563,s3287,s3294);
  not x1343(s3311,s3305);
  nand x1344(s2585,s3305,s3312);
  nand x1345(s2625,s3419,s3426);
  not x1346(s3283,s3277);
  nand x1347(s3286,s3277,s3284);
  nand x1348(s3304,s3295,s3302);
  not x1349(s3319,s3313);
  nand x1350(s3322,s3313,s3320);
  buf x1351(s3358,s2567);
  buf x1352(s3366,s2567);
  buf x1353(s3382,s2589);
  buf x1354(s3390,s2589);
  and x1355(s397,s330,s2514,s2657);
  and x1356(s2544,s330,s2508);
  nand x1357(s2562,s3290,s3293);
  nand x1358(s2584,s3308,s3311);
  not x1359(s3402,s3398);
  nand x1360(s2626,s2624,s2625);
  not x1361(s2632,s2629);
  and x1362(s2634,s2501,s2629);
  buf x1363(s2650,s2647);
  not x1364(s3268,s3264);
  buf x1365(s3256,s2508);
  nand x1366(s3285,s3280,s3283);
  nand x1367(s3321,s3316,s3319);
  nand x1368(s3371,s3303,s3304);
  buf x1369(s3403,s2609);
  buf x1370(s3411,s2609);
  or x1371(s362,s929,s933,s938);
  nor x1372(s1030,s929,s933,s938);
  or x1373(s399,s397,s398);
  nand x1374(s2564,s2562,s2563);
  not x1375(s3362,s3358);
  not x1376(s3370,s3366);
  nand x1377(s2586,s2584,s2585);
  not x1378(s3386,s3382);
  not x1379(s3394,s3390);
  and x1380(s2633,s330,s2505,s2632);
  buf x1381(s3261,s2527);
  buf x1382(s3269,s2527);
  nand x1383(s3347,s3285,s3286);
  nand x1384(s3395,s3321,s3322);
  not x1385(s363,s1030);
  nand x1386(s2536,s3256,s3259);
  not x1387(s3260,s3256);
  not x1388(s3377,s3371);
  nand x1389(s2580,s3371,s3378);
  not x1390(s3409,s3403);
  nand x1391(s2616,s3403,s3410);
  not x1392(s3417,s3411);
  nand x1393(s2622,s3411,s3418);
  nor x1394(s2635,s2633,s2634);
  and x1395(s2805,s2626,s2802);
  and x1396(s2808,s2626,s2803);
  buf x1397(s3334,s2544);
  buf x1398(s3342,s2544);
  buf x1399(s3454,s2650);
  and x1400(s364,s362,s363);
  nand x1401(s2537,s3253,s3260);
  not x1402(s3275,s3269);
  nand x1403(s2540,s3269,s3276);
  not x1404(s3353,s3347);
  nand x1405(s2557,s3347,s3354);
  nand x1406(s2579,s3374,s3377);
  not x1407(s3401,s3395);
  nand x1408(s2602,s3395,s3402);
  nand x1409(s2615,s3406,s3409);
  nand x1410(s2621,s3414,s3417);
  not x1411(s3267,s3261);
  nand x1412(s3112,s3261,s3268);
  buf x1413(s3355,s2564);
  buf x1414(s3363,s2564);
  buf x1415(s3379,s2586);
  buf x1416(s3387,s2586);
  nand x1417(s2538,s2536,s2537);
  nand x1418(s2539,s3272,s3275);
  not x1419(s3338,s3334);
  not x1420(s3346,s3342);
  nand x1421(s2556,s3350,s3353);
  nand x1422(s2581,s2579,s2580);
  nand x1423(s2601,s3398,s3401);
  nand x1424(s2617,s2615,s2616);
  nand x1425(s2623,s2621,s2622);
  buf x1426(s2638,s2635);
  not x1427(s3458,s3454);
  or x1428(s2814,s2805,s2808,s2811);
  nor x1429(s2816,s2805,s2808,s2811);
  nand x1430(s3111,s3264,s3267);
  nand x1431(s2541,s2539,s2540);
  nand x1432(s2558,s2556,s2557);
  not x1433(s3361,s3355);
  nand x1434(s2571,s3355,s3362);
  not x1435(s3369,s3363);
  nand x1436(s2577,s3363,s3370);
  not x1437(s3385,s3379);
  nand x1438(s2593,s3379,s3386);
  not x1439(s3393,s3387);
  nand x1440(s2598,s3387,s3394);
  nand x1441(s2603,s2601,s2602);
  nand x1442(s3113,s3111,s3112);
  and x1443(s3116,s330,s2538);
  not x1444(s3451,s2623);
  not x1445(s395,s2816);
  nand x1446(s2570,s3358,s3361);
  nand x1447(s2576,s3366,s3369);
  nand x1448(s2592,s3382,s3385);
  nand x1449(s2597,s3390,s3393);
  and x1450(s2736,s2581,s2733);
  and x1451(s2739,s2581,s2734);
  and x1452(s2788,s2617,s2785);
  buf x1453(s3438,s2638);
  and x1454(s3446,s2617,s2647);
  buf x1455(s3459,s2814);
  and x1456(s396,s2814,s395);
  not x1457(s3119,s3113);
  not x1458(s3120,s3116);
  nand x1459(s2572,s2570,s2571);
  nand x1460(s2578,s2576,s2577);
  nand x1461(s2594,s2592,s2593);
  nand x1462(s2599,s2597,s2598);
  nand x1463(s2677,s3451,s3458);
  not x1464(s3457,s3451);
  and x1465(s2700,s2558,s2697);
  and x1466(s2771,s2603,s2768);
  buf x1467(s3331,s2541);
  buf x1468(s3339,s2541);
  buf x1469(s3427,s2558);
  buf x1470(s3443,s2603);
  nand x1471(s954,s3116,s3119);
  nand x1472(s955,s3113,s3120);
  not x1473(s2600,s2599);
  not x1474(s3442,s3438);
  not x1475(s3450,s3446);
  nand x1476(s2676,s3454,s3457);
  or x1477(s2745,s2736,s2739,s2742);
  nor x1478(s2748,s2736,s2739,s2742);
  not x1479(s3465,s3459);
  not x1480(s3435,s2578);
  nand x1481(s950,s954,s955);
  not x1482(s3337,s3331);
  nand x1483(s2548,s3331,s3338);
  not x1484(s3345,s3339);
  nand x1485(s2553,s3339,s3346);
  nor x1486(s2661,s2600,s2650);
  and x1487(s2662,s2617,s2603,s2594,s2650);
  not x1488(s3433,s3427);
  not x1489(s3449,s3443);
  nand x1490(s2672,s3443,s3450);
  nand x1491(s2674,s2676,s2677);
  and x1492(s2719,s2572,s2716);
  and x1493(s2754,s2594,s2751);
  and x1494(s3430,s2572,s2635);
  not x1495(s383,s2748);
  and x1496(s951,s950,s943);
  nand x1497(s2547,s3334,s3337);
  nand x1498(s2552,s3342,s3345);
  or x1499(s2663,s2661,s2662);
  nand x1500(s2670,s3435,s3442);
  not x1501(s3441,s3435);
  nand x1502(s2671,s3446,s3449);
  not x1503(s2675,s2674);
  buf x1504(s3491,s2745);
  buf x1505(s3499,s2745);
  and x1506(s384,s2745,s383);
  nand x1507(s2549,s2547,s2548);
  nand x1508(s2554,s2552,s2553);
  nand x1509(s2664,s3430,s3433);
  not x1510(s3434,s3430);
  nand x1511(s2669,s3438,s3441);
  nand x1512(s2673,s2671,s2672);
  and x1513(s2757,s2663,s2752);
  and x1514(s2791,s2675,s2786);
  or x1515(s365,s944,s947,s951);
  nor x1516(s1031,s944,s947,s951);
  not x1517(s2555,s2554);
  nand x1518(s2665,s3427,s3434);
  nand x1519(s2667,s2669,s2670);
  and x1520(s2774,s2673,s2769);
  not x1521(s3497,s3491);
  not x1522(s3505,s3499);
  not x1523(s366,s1031);
  nor x1524(s2658,s2555,s2638);
  and x1525(s2659,s2572,s2558,s2549,s2638);
  nand x1526(s2666,s2664,s2665);
  not x1527(s2668,s2667);
  and x1528(s2681,s2549,s2678);
  or x1529(s2763,s2754,s2757,s2760);
  nor x1530(s2765,s2754,s2757,s2760);
  or x1531(s2797,s2788,s2791,s2794);
  nor x1532(s2799,s2788,s2791,s2794);
  and x1533(s367,s365,s366);
  or x1534(s2660,s2658,s2659);
  and x1535(s2703,s2666,s2698);
  and x1536(s2722,s2668,s2717);
  or x1537(s2780,s2771,s2774,s2777);
  nor x1538(s2782,s2771,s2774,s2777);
  not x1539(s386,s2765);
  not x1540(s392,s2799);
  and x1541(s2684,s2660,s2679);
  buf x1542(s3462,s2797);
  buf x1543(s3470,s2763);
  and x1544(s387,s2763,s386);
  not x1545(s389,s2782);
  and x1546(s393,s2797,s392);
  or x1547(s2709,s2700,s2703,s2706);
  nor x1548(s2713,s2700,s2703,s2706);
  or x1549(s2728,s2719,s2722,s2725);
  nor x1550(s2730,s2719,s2722,s2725);
  and x1551(s2922,s2816,s2799,s2782,s2765);
  buf x1552(s3467,s2780);
  and x1553(s390,s2780,s389);
  or x1554(s2690,s2681,s2684,s2687);
  nor x1555(s2694,s2681,s2684,s2687);
  nand x1556(s2821,s3462,s3465);
  not x1557(s3466,s3462);
  not x1558(s3474,s3470);
  and x1559(s378,s2709,s2709);
  not x1560(s380,s2730);
  nand x1561(s2822,s3459,s3466);
  not x1562(s3473,s3467);
  nand x1563(s2827,s3467,s3474);
  buf x1564(s2839,s2728);
  and x1565(s2883,s2709,s2871);
  buf x1566(s3507,s2709);
  and x1567(s375,s2690,s2690);
  and x1568(s381,s2728,s380);
  nand x1569(s2823,s2821,s2822);
  nand x1570(s2826,s3470,s3473);
  and x1571(s2880,s2871,s2690);
  and x1572(s2925,s2748,s2730,s2713,s2694);
  and x1573(s2928,s2713,s2694,s2874);
  buf x1574(s3510,s2690);
  nand x1575(s2828,s2826,s2827);
  buf x1576(s3494,s2839);
  buf x1577(s3502,s2839);
  not x1578(s3513,s3507);
  buf x1579(s3544,s2883);
  buf x1580(s3552,s2883);
  and x1581(s406,s2922,s2925);
  and x1582(s2929,s2922,s2925);
  buf x1583(s3475,s2823);
  buf x1584(s3483,s2823);
  not x1585(s3514,s3510);
  nand x1586(s3515,s3510,s3513);
  buf x1587(s3541,s2880);
  buf x1588(s3549,s2880);
  not x1589(s407,s406);
  nor x1590(s2930,s2928,s2929);
  nand x1591(s2842,s3494,s3497);
  not x1592(s3498,s3494);
  nand x1593(s2852,s3502,s3505);
  not x1594(s3506,s3502);
  not x1595(s3548,s3544);
  not x1596(s3556,s3552);
  buf x1597(s3478,s2828);
  buf x1598(s3486,s2828);
  nand x1599(s3516,s3507,s3514);
  and x1600(s408,s213,s2930);
  not x1601(s3481,s3475);
  not x1602(s3489,s3483);
  nand x1603(s2843,s3491,s3498);
  nand x1604(s2853,s3499,s3506);
  not x1605(s3547,s3541);
  nand x1606(s2887,s3541,s3548);
  nand x1607(s2896,s3549,s3556);
  not x1608(s3555,s3549);
  nand x1609(s3520,s3515,s3516);
  not x1610(s409,s408);
  nand x1611(s2831,s3478,s3481);
  not x1612(s3482,s3478);
  nand x1613(s2836,s3486,s3489);
  not x1614(s3490,s3486);
  nand x1615(s2844,s2842,s2843);
  nand x1616(s2848,s2852,s2853);
  nand x1617(s2886,s3544,s3547);
  nand x1618(s2895,s3552,s3555);
  nand x1619(s2832,s3475,s3482);
  nand x1620(s2837,s3483,s3490);
  not x1621(s2849,s2848);
  not x1622(s3524,s3520);
  nand x1623(s2888,s2886,s2887);
  nand x1624(s2891,s2895,s2896);
  nand x1625(s2833,s2831,s2832);
  nand x1626(s2838,s2836,s2837);
  not x1627(s2892,s2891);
  buf x1628(s3517,s2844);
  and x1629(s2906,s2844,s2888,s2900);
  and x1630(s2908,s2849,s2888,s2903);
  not x1631(s2913,s2838);
  not x1632(s3523,s3517);
  nand x1633(s2855,s3517,s3524);
  and x1634(s2907,s2844,s2892,s2903);
  and x1635(s2909,s2849,s2892,s2900);
  buf x1636(s3525,s2833);
  buf x1637(s3533,s2833);
  nand x1638(s2854,s3520,s3523);
  or x1639(s2910,s2906,s2907,s2908,s2909);
  buf x1640(s3560,s2913);
  buf x1641(s3568,s2913);
  nand x1642(s2856,s2854,s2855);
  not x1643(s3539,s3533);
  not x1644(s3531,s3525);
  not x1645(s3572,s3568);
  not x1646(s3564,s3560);
  buf x1647(s3557,s2910);
  buf x1648(s3565,s2910);
  buf x1649(s3528,s2856);
  buf x1650(s3536,s2856);
  nand x1651(s2921,s3557,s3564);
  nand x1652(s2917,s3565,s3572);
  not x1653(s3571,s3565);
  not x1654(s3563,s3557);
  nand x1655(s2863,s3528,s3531);
  nand x1656(s2859,s3536,s3539);
  nand x1657(s2920,s3560,s3563);
  nand x1658(s2916,s3568,s3571);
  not x1659(s3540,s3536);
  not x1660(s3532,s3528);
  nand x1661(s2864,s3525,s3532);
  nand x1662(s2860,s3533,s3540);
  nand x1663(s403,s2920,s2921);
  nand x1664(s404,s2916,s2917);
  nand x1665(s400,s2863,s2864);
  nand x1666(s401,s2859,s2860);
  and x1667(s405,s403,s404);
  nand x1668(s402,s400,s401);

endmodule
