module c432(s223gat,s329gat,s370gat,s421gat,s430gat,s431gat,s432gat,s1gat,s4gat,s8gat,s11gat,s14gat,s17gat,s21gat,s24gat,s27gat,s30gat,s34gat,s37gat,s40gat,s43gat,s47gat,s50gat,s53gat,s56gat,s60gat,s63gat,s66gat,s69gat,s73gat,s76gat,s79gat,s82gat,s86gat,s89gat,s92gat,s95gat,s99gat,s102gat,s105gat,s108gat,s112gat,s115gat);

  output s223gat;
  output s329gat;
  output s370gat;
  output s421gat;
  output s430gat;
  output s431gat;
  output s432gat;
  input s1gat;
  input s4gat;
  input s8gat;
  input s11gat;
  input s14gat;
  input s17gat;
  input s21gat;
  input s24gat;
  input s27gat;
  input s30gat;
  input s34gat;
  input s37gat;
  input s40gat;
  input s43gat;
  input s47gat;
  input s50gat;
  input s53gat;
  input s56gat;
  input s60gat;
  input s63gat;
  input s66gat;
  input s69gat;
  input s73gat;
  input s76gat;
  input s79gat;
  input s82gat;
  input s86gat;
  input s89gat;
  input s92gat;
  input s95gat;
  input s99gat;
  input s102gat;
  input s105gat;
  input s108gat;
  input s112gat;
  input s115gat;

  not x0(s118gat,s1gat);
  not x1(s119gat,s4gat);
  not x2(s122gat,s11gat);
  not x3(s123gat,s17gat);
  not x4(s126gat,s24gat);
  not x5(s127gat,s30gat);
  not x6(s130gat,s37gat);
  not x7(s131gat,s43gat);
  not x8(s134gat,s50gat);
  not x9(s135gat,s56gat);
  not x10(s138gat,s63gat);
  not x11(s139gat,s69gat);
  not x12(s142gat,s76gat);
  not x13(s143gat,s82gat);
  not x14(s146gat,s89gat);
  not x15(s147gat,s95gat);
  not x16(s150gat,s102gat);
  not x17(s151gat,s108gat);
  nand x18(s154gat,s118gat,s4gat);
  nor x19(s157gat,s8gat,s119gat);
  nor x20(s158gat,s14gat,s119gat);
  nand x21(s159gat,s122gat,s17gat);
  nand x22(s162gat,s126gat,s30gat);
  nand x23(s165gat,s130gat,s43gat);
  nand x24(s168gat,s134gat,s56gat);
  nand x25(s171gat,s138gat,s69gat);
  nand x26(s174gat,s142gat,s82gat);
  nand x27(s177gat,s146gat,s95gat);
  nand x28(s180gat,s150gat,s108gat);
  nor x29(s183gat,s21gat,s123gat);
  nor x30(s184gat,s27gat,s123gat);
  nor x31(s185gat,s34gat,s127gat);
  nor x32(s186gat,s40gat,s127gat);
  nor x33(s187gat,s47gat,s131gat);
  nor x34(s188gat,s53gat,s131gat);
  nor x35(s189gat,s60gat,s135gat);
  nor x36(s190gat,s66gat,s135gat);
  nor x37(s191gat,s73gat,s139gat);
  nor x38(s192gat,s79gat,s139gat);
  nor x39(s193gat,s86gat,s143gat);
  nor x40(s194gat,s92gat,s143gat);
  nor x41(s195gat,s99gat,s147gat);
  nor x42(s196gat,s105gat,s147gat);
  nor x43(s197gat,s112gat,s151gat);
  nor x44(s198gat,s115gat,s151gat);
  and x45(s199gat,s154gat,s159gat,s162gat,s165gat,s168gat,s171gat,s174gat,s177gat,s180gat);
  not x46(s203gat,s199gat);
  not x47(s213gat,s199gat);
  not x48(s223gat,s199gat);
  xor x49(s224gat,s203gat,s154gat);
  xor x50(s227gat,s203gat,s159gat);
  xor x51(s230gat,s203gat,s162gat);
  xor x52(s233gat,s203gat,s165gat);
  xor x53(s236gat,s203gat,s168gat);
  xor x54(s239gat,s203gat,s171gat);
  nand x55(s242gat,s1gat,s213gat);
  xor x56(s243gat,s203gat,s174gat);
  nand x57(s246gat,s213gat,s11gat);
  xor x58(s247gat,s203gat,s177gat);
  nand x59(s250gat,s213gat,s24gat);
  xor x60(s251gat,s203gat,s180gat);
  nand x61(s254gat,s213gat,s37gat);
  nand x62(s255gat,s213gat,s50gat);
  nand x63(s256gat,s213gat,s63gat);
  nand x64(s257gat,s213gat,s76gat);
  nand x65(s258gat,s213gat,s89gat);
  nand x66(s259gat,s213gat,s102gat);
  nand x67(s260gat,s224gat,s157gat);
  nand x68(s263gat,s224gat,s158gat);
  nand x69(s264gat,s227gat,s183gat);
  nand x70(s267gat,s230gat,s185gat);
  nand x71(s270gat,s233gat,s187gat);
  nand x72(s273gat,s236gat,s189gat);
  nand x73(s276gat,s239gat,s191gat);
  nand x74(s279gat,s243gat,s193gat);
  nand x75(s282gat,s247gat,s195gat);
  nand x76(s285gat,s251gat,s197gat);
  nand x77(s288gat,s227gat,s184gat);
  nand x78(s289gat,s230gat,s186gat);
  nand x79(s290gat,s233gat,s188gat);
  nand x80(s291gat,s236gat,s190gat);
  nand x81(s292gat,s239gat,s192gat);
  nand x82(s293gat,s243gat,s194gat);
  nand x83(s294gat,s247gat,s196gat);
  nand x84(s295gat,s251gat,s198gat);
  and x85(s296gat,s260gat,s264gat,s267gat,s270gat,s273gat,s276gat,s279gat,s282gat,s285gat);
  not x86(s300gat,s263gat);
  not x87(s301gat,s288gat);
  not x88(s302gat,s289gat);
  not x89(s303gat,s290gat);
  not x90(s304gat,s291gat);
  not x91(s305gat,s292gat);
  not x92(s306gat,s293gat);
  not x93(s307gat,s294gat);
  not x94(s308gat,s295gat);
  not x95(s309gat,s296gat);
  not x96(s319gat,s296gat);
  not x97(s329gat,s296gat);
  xor x98(s330gat,s309gat,s260gat);
  xor x99(s331gat,s309gat,s264gat);
  xor x100(s332gat,s309gat,s267gat);
  xor x101(s333gat,s309gat,s270gat);
  nand x102(s334gat,s8gat,s319gat);
  xor x103(s335gat,s309gat,s273gat);
  nand x104(s336gat,s319gat,s21gat);
  xor x105(s337gat,s309gat,s276gat);
  nand x106(s338gat,s319gat,s34gat);
  xor x107(s339gat,s309gat,s279gat);
  nand x108(s340gat,s319gat,s47gat);
  xor x109(s341gat,s309gat,s282gat);
  nand x110(s342gat,s319gat,s60gat);
  xor x111(s343gat,s309gat,s285gat);
  nand x112(s344gat,s319gat,s73gat);
  nand x113(s345gat,s319gat,s86gat);
  nand x114(s346gat,s319gat,s99gat);
  nand x115(s347gat,s319gat,s112gat);
  nand x116(s348gat,s330gat,s300gat);
  nand x117(s349gat,s331gat,s301gat);
  nand x118(s350gat,s332gat,s302gat);
  nand x119(s351gat,s333gat,s303gat);
  nand x120(s352gat,s335gat,s304gat);
  nand x121(s353gat,s337gat,s305gat);
  nand x122(s354gat,s339gat,s306gat);
  nand x123(s355gat,s341gat,s307gat);
  nand x124(s356gat,s343gat,s308gat);
  and x125(s357gat,s348gat,s349gat,s350gat,s351gat,s352gat,s353gat,s354gat,s355gat,s356gat);
  not x126(s360gat,s357gat);
  not x127(s370gat,s357gat);
  nand x128(s371gat,s14gat,s360gat);
  nand x129(s372gat,s360gat,s27gat);
  nand x130(s373gat,s360gat,s40gat);
  nand x131(s374gat,s360gat,s53gat);
  nand x132(s375gat,s360gat,s66gat);
  nand x133(s376gat,s360gat,s79gat);
  nand x134(s377gat,s360gat,s92gat);
  nand x135(s378gat,s360gat,s105gat);
  nand x136(s379gat,s360gat,s115gat);
  nand x137(s380gat,s4gat,s242gat,s334gat,s371gat);
  nand x138(s381gat,s246gat,s336gat,s372gat,s17gat);
  nand x139(s386gat,s250gat,s338gat,s373gat,s30gat);
  nand x140(s393gat,s254gat,s340gat,s374gat,s43gat);
  nand x141(s399gat,s255gat,s342gat,s375gat,s56gat);
  nand x142(s404gat,s256gat,s344gat,s376gat,s69gat);
  nand x143(s407gat,s257gat,s345gat,s377gat,s82gat);
  nand x144(s411gat,s258gat,s346gat,s378gat,s95gat);
  nand x145(s414gat,s259gat,s347gat,s379gat,s108gat);
  not x146(s415gat,s380gat);
  and x147(s416gat,s381gat,s386gat,s393gat,s399gat,s404gat,s407gat,s411gat,s414gat);
  not x148(s417gat,s393gat);
  not x149(s418gat,s404gat);
  not x150(s419gat,s407gat);
  not x151(s420gat,s411gat);
  nor x152(s421gat,s415gat,s416gat);
  nand x153(s422gat,s386gat,s417gat);
  nand x154(s425gat,s386gat,s393gat,s418gat,s399gat);
  nand x155(s428gat,s399gat,s393gat,s419gat);
  nand x156(s429gat,s386gat,s393gat,s407gat,s420gat);
  nand x157(s430gat,s381gat,s386gat,s422gat,s399gat);
  nand x158(s431gat,s381gat,s386gat,s425gat,s428gat);
  nand x159(s432gat,s381gat,s422gat,s425gat,s429gat);

endmodule
