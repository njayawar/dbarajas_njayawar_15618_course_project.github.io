module c5315(s144,s298,s973,s594,s599,s600,s601,s602,s603,s604,s611,s612,s810,s848,s849,s850,s851,s634,s815,s845,s847,s926,s923,s921,s892,s887,s606,s656,s809,s993,s978,s949,s939,s889,s593,s636,s704,s717,s820,s639,s673,s707,s715,s598,s610,s588,s615,s626,s632,s1002,s1004,s591,s618,s621,s629,s822,s838,s861,s623,s722,s832,s834,s836,s859,s871,s873,s875,s877,s998,s1000,s575,s585,s661,s693,s747,s752,s757,s762,s787,s792,s797,s802,s642,s664,s667,s670,s676,s696,s699,s702,s818,s813,s824,s826,s828,s830,s854,s863,s865,s867,s869,s712,s727,s732,s737,s742,s772,s777,s782,s645,s648,s651,s654,s679,s682,s685,s688,s843,s882,s767,s807,s658,s690,s1,s4,s11,s14,s17,s20,s23,s24,s25,s26,s27,s31,s34,s37,s40,s43,s46,s49,s52,s53,s54,s61,s64,s67,s70,s73,s76,s79,s80,s81,s82,s83,s86,s87,s88,s91,s94,s97,s100,s103,s106,s109,s112,s113,s114,s115,s116,s117,s118,s119,s120,s121,s122,s123,s126,s127,s128,s129,s130,s131,s132,s135,s136,s137,s140,s141,s145,s146,s149,s152,s155,s158,s161,s164,s167,s170,s173,s176,s179,s182,s185,s188,s191,s194,s197,s200,s203,s206,s209,s210,s217,s218,s225,s226,s233,s234,s241,s242,s245,s248,s251,s254,s257,s264,s265,s272,s273,s280,s281,s288,s289,s292,s293,s299,s302,s307,s308,s315,s316,s323,s324,s331,s332,s335,s338,s341,s348,s351,s358,s361,s366,s369,s372,s373,s374,s386,s389,s400,s411,s422,s435,s446,s457,s468,s479,s490,s503,s514,s523,s534,s545,s549,s552,s556,s559,s562,s1497,s1689,s1690,s1691,s1694,s2174,s2358,s2824,s3173,s3546,s3548,s3550,s3552,s3717,s3724,s4087,s4088,s4089,s4090,s4091,s4092,s4115);

  output s144;
  output s298;
  output s973;
  output s594;
  output s599;
  output s600;
  output s601;
  output s602;
  output s603;
  output s604;
  output s611;
  output s612;
  output s810;
  output s848;
  output s849;
  output s850;
  output s851;
  output s634;
  output s815;
  output s845;
  output s847;
  output s926;
  output s923;
  output s921;
  output s892;
  output s887;
  output s606;
  output s656;
  output s809;
  output s993;
  output s978;
  output s949;
  output s939;
  output s889;
  output s593;
  output s636;
  output s704;
  output s717;
  output s820;
  output s639;
  output s673;
  output s707;
  output s715;
  output s598;
  output s610;
  output s588;
  output s615;
  output s626;
  output s632;
  output s1002;
  output s1004;
  output s591;
  output s618;
  output s621;
  output s629;
  output s822;
  output s838;
  output s861;
  output s623;
  output s722;
  output s832;
  output s834;
  output s836;
  output s859;
  output s871;
  output s873;
  output s875;
  output s877;
  output s998;
  output s1000;
  output s575;
  output s585;
  output s661;
  output s693;
  output s747;
  output s752;
  output s757;
  output s762;
  output s787;
  output s792;
  output s797;
  output s802;
  output s642;
  output s664;
  output s667;
  output s670;
  output s676;
  output s696;
  output s699;
  output s702;
  output s818;
  output s813;
  output s824;
  output s826;
  output s828;
  output s830;
  output s854;
  output s863;
  output s865;
  output s867;
  output s869;
  output s712;
  output s727;
  output s732;
  output s737;
  output s742;
  output s772;
  output s777;
  output s782;
  output s645;
  output s648;
  output s651;
  output s654;
  output s679;
  output s682;
  output s685;
  output s688;
  output s843;
  output s882;
  output s767;
  output s807;
  output s658;
  output s690;
  input s1;
  input s4;
  input s11;
  input s14;
  input s17;
  input s20;
  input s23;
  input s24;
  input s25;
  input s26;
  input s27;
  input s31;
  input s34;
  input s37;
  input s40;
  input s43;
  input s46;
  input s49;
  input s52;
  input s53;
  input s54;
  input s61;
  input s64;
  input s67;
  input s70;
  input s73;
  input s76;
  input s79;
  input s80;
  input s81;
  input s82;
  input s83;
  input s86;
  input s87;
  input s88;
  input s91;
  input s94;
  input s97;
  input s100;
  input s103;
  input s106;
  input s109;
  input s112;
  input s113;
  input s114;
  input s115;
  input s116;
  input s117;
  input s118;
  input s119;
  input s120;
  input s121;
  input s122;
  input s123;
  input s126;
  input s127;
  input s128;
  input s129;
  input s130;
  input s131;
  input s132;
  input s135;
  input s136;
  input s137;
  input s140;
  input s141;
  input s145;
  input s146;
  input s149;
  input s152;
  input s155;
  input s158;
  input s161;
  input s164;
  input s167;
  input s170;
  input s173;
  input s176;
  input s179;
  input s182;
  input s185;
  input s188;
  input s191;
  input s194;
  input s197;
  input s200;
  input s203;
  input s206;
  input s209;
  input s210;
  input s217;
  input s218;
  input s225;
  input s226;
  input s233;
  input s234;
  input s241;
  input s242;
  input s245;
  input s248;
  input s251;
  input s254;
  input s257;
  input s264;
  input s265;
  input s272;
  input s273;
  input s280;
  input s281;
  input s288;
  input s289;
  input s292;
  input s293;
  input s299;
  input s302;
  input s307;
  input s308;
  input s315;
  input s316;
  input s323;
  input s324;
  input s331;
  input s332;
  input s335;
  input s338;
  input s341;
  input s348;
  input s351;
  input s358;
  input s361;
  input s366;
  input s369;
  input s372;
  input s373;
  input s374;
  input s386;
  input s389;
  input s400;
  input s411;
  input s422;
  input s435;
  input s446;
  input s457;
  input s468;
  input s479;
  input s490;
  input s503;
  input s514;
  input s523;
  input s534;
  input s545;
  input s549;
  input s552;
  input s556;
  input s559;
  input s562;
  input s1497;
  input s1689;
  input s1690;
  input s1691;
  input s1694;
  input s2174;
  input s2358;
  input s2824;
  input s3173;
  input s3546;
  input s3548;
  input s3550;
  input s3552;
  input s3717;
  input s3724;
  input s4087;
  input s4088;
  input s4089;
  input s4090;
  input s4091;
  input s4092;
  input s4115;

  buf x0(s144,s141);
  buf x1(s298,s293);
  and x2(s4114,s135,s4115);
  not x3(s2825,s2824);
  buf x4(s973,s3173);
  not x5(s3547,s3546);
  not x6(s3549,s3548);
  not x7(s3551,s3550);
  not x8(s3553,s3552);
  not x9(s594,s545);
  not x10(s599,s348);
  not x11(s600,s366);
  and x12(s601,s552,s562);
  not x13(s602,s549);
  not x14(s603,s545);
  not x15(s604,s545);
  not x16(s611,s338);
  not x17(s612,s358);
  nand x18(s633,s373,s1);
  and x19(s810,s141,s145);
  not x20(s814,s3173);
  not x21(s816,s4114);
  and x22(s844,s2825,s27);
  and x23(s846,s386,s556);
  not x24(s848,s245);
  not x25(s849,s552);
  not x26(s850,s562);
  not x27(s851,s559);
  and x28(s852,s386,s559,s556,s552);
  not x29(s1502,s1497);
  buf x30(s1528,s1689);
  buf x31(s1552,s1690);
  buf x32(s1609,s1689);
  buf x33(s1633,s1690);
  buf x34(s1697,s137);
  buf x35(s1698,s137);
  buf x36(s1701,s141);
  not x37(s2179,s2174);
  buf x38(s2203,s1691);
  buf x39(s2226,s1694);
  buf x40(s2281,s1691);
  buf x41(s2304,s1694);
  buf x42(s2361,s254);
  buf x43(s2370,s251);
  buf x44(s2382,s251);
  buf x45(s2393,s248);
  buf x46(s2405,s248);
  buf x47(s2418,s4088);
  buf x48(s2442,s4087);
  buf x49(s2476,s4089);
  buf x50(s2500,s4090);
  buf x51(s2533,s210);
  buf x52(s2537,s210);
  buf x53(s2541,s218);
  buf x54(s2545,s218);
  buf x55(s2549,s226);
  buf x56(s2553,s226);
  buf x57(s2557,s234);
  buf x58(s2561,s234);
  buf x59(s2627,s257);
  buf x60(s2631,s257);
  buf x61(s2635,s265);
  buf x62(s2639,s265);
  buf x63(s2643,s273);
  buf x64(s2647,s273);
  buf x65(s2651,s281);
  buf x66(s2655,s281);
  buf x67(s2721,s335);
  buf x68(s2734,s335);
  buf x69(s2816,s206);
  and x70(s2822,s27,s31);
  buf x71(s2826,s1);
  buf x72(s2828,s2358);
  buf x73(s2882,s293);
  buf x74(s2886,s302);
  buf x75(s2890,s308);
  buf x76(s2894,s308);
  buf x77(s2898,s316);
  buf x78(s2902,s316);
  buf x79(s2948,s324);
  buf x80(s2952,s324);
  buf x81(s2956,s341);
  buf x82(s2960,s341);
  buf x83(s2964,s351);
  buf x84(s2968,s351);
  buf x85(s3024,s257);
  buf x86(s3028,s257);
  buf x87(s3032,s265);
  buf x88(s3036,s265);
  buf x89(s3040,s273);
  buf x90(s3044,s273);
  buf x91(s3048,s281);
  buf x92(s3052,s281);
  buf x93(s3092,s332);
  buf x94(s3105,s332);
  buf x95(s3175,s549);
  and x96(s3176,s31,s27);
  not x97(s3181,s2358);
  buf x98(s3204,s324);
  buf x99(s3208,s324);
  buf x100(s3212,s341);
  buf x101(s3216,s341);
  buf x102(s3220,s351);
  buf x103(s3224,s351);
  buf x104(s3256,s293);
  buf x105(s3260,s302);
  buf x106(s3264,s308);
  buf x107(s3268,s308);
  buf x108(s3272,s316);
  buf x109(s3276,s316);
  buf x110(s3302,s361);
  buf x111(s3314,s361);
  buf x112(s3354,s210);
  buf x113(s3358,s210);
  buf x114(s3362,s218);
  buf x115(s3366,s218);
  buf x116(s3370,s226);
  buf x117(s3374,s226);
  buf x118(s3378,s234);
  buf x119(s3382,s234);
  not x120(s3440,s324);
  buf x121(s3554,s242);
  buf x122(s3555,s242);
  buf x123(s3556,s254);
  buf x124(s3558,s4088);
  buf x125(s3582,s4087);
  buf x126(s3616,s4092);
  buf x127(s3628,s4091);
  buf x128(s3660,s4089);
  buf x129(s3684,s4090);
  not x130(s3721,s3717);
  not x131(s3728,s3724);
  buf x132(s3737,s4091);
  buf x133(s3757,s4092);
  buf x134(s3795,s4091);
  buf x135(s3815,s4092);
  buf x136(s3972,s4091);
  buf x137(s3991,s4092);
  buf x138(s4030,s4091);
  buf x139(s4049,s4092);
  buf x140(s4110,s299);
  buf x141(s4119,s446);
  buf x142(s4127,s457);
  buf x143(s4135,s468);
  buf x144(s4143,s422);
  buf x145(s4151,s435);
  buf x146(s4159,s389);
  buf x147(s4167,s400);
  buf x148(s4175,s411);
  buf x149(s4183,s374);
  buf x150(s4188,s4);
  buf x151(s4276,s446);
  buf x152(s4284,s457);
  buf x153(s4292,s468);
  buf x154(s4300,s435);
  buf x155(s4308,s389);
  buf x156(s4316,s400);
  buf x157(s4324,s411);
  buf x158(s4332,s422);
  buf x159(s4340,s374);
  buf x160(s4631,s479);
  buf x161(s4639,s490);
  buf x162(s4647,s503);
  buf x163(s4655,s514);
  buf x164(s4663,s523);
  buf x165(s4671,s534);
  buf x166(s4676,s54);
  buf x167(s4764,s479);
  buf x168(s4772,s503);
  buf x169(s4780,s514);
  buf x170(s4788,s523);
  buf x171(s4796,s534);
  buf x172(s4804,s490);
  buf x173(s5082,s361);
  buf x174(s5085,s369);
  buf x175(s5090,s341);
  buf x176(s5093,s351);
  buf x177(s5098,s308);
  buf x178(s5101,s316);
  buf x179(s5108,s293);
  buf x180(s5111,s302);
  buf x181(s5332,s281);
  buf x182(s5335,s289);
  buf x183(s5340,s265);
  buf x184(s5343,s273);
  buf x185(s5348,s234);
  buf x186(s5351,s257);
  buf x187(s5356,s218);
  buf x188(s5359,s226);
  buf x189(s5369,s210);
  not x190(s634,s633);
  and x191(s815,s136,s814);
  not x192(s845,s844);
  not x193(s847,s846);
  buf x194(s926,s1697);
  buf x195(s923,s1701);
  buf x196(s921,s2826);
  and x197(s2979,s3553,s514);
  or x198(s2999,s3547,s514);
  buf x199(s892,s3175);
  buf x200(s887,s4110);
  not x201(s606,s3175);
  and x202(s1580,s170,s1528,s1552);
  and x203(s1586,s173,s1528,s1552);
  and x204(s1592,s167,s1528,s1552);
  and x205(s1598,s164,s1528,s1552);
  and x206(s1604,s161,s1528,s1552);
  nand x207(s656,s2822,s140);
  and x208(s1668,s185,s1609,s1633);
  and x209(s1674,s158,s1609,s1633);
  and x210(s1680,s152,s1609,s1633);
  and x211(s1686,s146,s1609,s1633);
  and x212(s2254,s170,s2203,s2226);
  and x213(s2260,s173,s2203,s2226);
  and x214(s2266,s167,s2203,s2226);
  and x215(s2272,s164,s2203,s2226);
  and x216(s2278,s161,s2203,s2226);
  and x217(s2339,s185,s2281,s2304);
  and x218(s2345,s158,s2281,s2304);
  and x219(s2351,s152,s2281,s2304);
  and x220(s2357,s146,s2281,s2304);
  and x221(s711,s106,s3660,s3684);
  and x222(s721,s61,s2418,s2442);
  and x223(s726,s106,s3558,s3582);
  and x224(s731,s49,s3558,s3582);
  and x225(s736,s103,s3558,s3582);
  and x226(s741,s40,s3558,s3582);
  and x227(s746,s37,s3558,s3582);
  and x228(s751,s20,s2418,s2442);
  and x229(s756,s17,s2418,s2442);
  and x230(s761,s70,s2418,s2442);
  and x231(s766,s64,s2418,s2442);
  and x232(s771,s49,s3660,s3684);
  and x233(s776,s103,s3660,s3684);
  and x234(s781,s40,s3660,s3684);
  and x235(s786,s37,s3660,s3684);
  and x236(s791,s20,s2476,s2500);
  and x237(s796,s17,s2476,s2500);
  and x238(s801,s70,s2476,s2500);
  and x239(s806,s64,s2476,s2500);
  not x240(s809,s2822);
  and x241(s3734,s123,s3728,s3717);
  and x242(s842,s3795,s3815);
  and x243(s858,s61,s2476,s2500);
  and x244(s881,s3737,s3757);
  not x245(s4123,s4119);
  not x246(s4131,s4127);
  not x247(s4139,s4135);
  not x248(s4147,s4143);
  not x249(s4155,s4151);
  not x250(s4163,s4159);
  not x251(s4171,s4167);
  not x252(s4179,s4175);
  not x253(s4187,s4183);
  not x254(s4194,s4188);
  not x255(s4282,s4276);
  not x256(s4290,s4284);
  not x257(s4298,s4292);
  not x258(s4306,s4300);
  not x259(s4314,s4308);
  not x260(s4322,s4316);
  not x261(s4330,s4324);
  not x262(s4338,s4332);
  not x263(s4346,s4340);
  buf x264(s1526,s1697);
  not x265(s1540,s1528);
  not x266(s1564,s1552);
  buf x267(s1606,s1697);
  not x268(s1621,s1609);
  not x269(s1645,s1633);
  and x270(s1661,s179,s1609,s1633);
  buf x271(s1688,s2826);
  not x272(s4635,s4631);
  not x273(s4643,s4639);
  not x274(s4651,s4647);
  not x275(s4659,s4655);
  not x276(s4667,s4663);
  not x277(s4675,s4671);
  not x278(s4682,s4676);
  not x279(s4770,s4764);
  not x280(s4778,s4772);
  not x281(s4786,s4780);
  not x282(s4794,s4788);
  not x283(s4802,s4796);
  not x284(s4810,s4804);
  buf x285(s2202,s1698);
  not x286(s2215,s2203);
  not x287(s2238,s2226);
  buf x288(s2279,s1698);
  not x289(s2293,s2281);
  not x290(s2316,s2304);
  and x291(s2332,s179,s2281,s2304);
  not x292(s2430,s2418);
  not x293(s2454,s2442);
  not x294(s2488,s2476);
  not x295(s2512,s2500);
  not x296(s2536,s2533);
  not x297(s2540,s2537);
  not x298(s2544,s2541);
  not x299(s2548,s2545);
  not x300(s2552,s2549);
  not x301(s2556,s2553);
  not x302(s2560,s2557);
  not x303(s2564,s2561);
  and x304(s2566,s3553,s457,s2537);
  and x305(s2572,s3553,s468,s2545);
  and x306(s2578,s3553,s422,s2553);
  and x307(s2584,s3553,s435,s2561);
  and x308(s2590,s3547,s2533);
  and x309(s2595,s3547,s2541);
  and x310(s2600,s3547,s2549);
  and x311(s2605,s3547,s2557);
  not x312(s2630,s2627);
  not x313(s2634,s2631);
  not x314(s2638,s2635);
  not x315(s2642,s2639);
  not x316(s2646,s2643);
  not x317(s2650,s2647);
  not x318(s2654,s2651);
  not x319(s2658,s2655);
  and x320(s2660,s3553,s389,s2631);
  and x321(s2666,s3553,s400,s2639);
  and x322(s2672,s3553,s411,s2647);
  and x323(s2678,s3553,s374,s2655);
  and x324(s2684,s3547,s2627);
  and x325(s2689,s3547,s2635);
  and x326(s2694,s3547,s2643);
  and x327(s2699,s3547,s2651);
  not x328(s2728,s2721);
  not x329(s2741,s2734);
  and x330(s2748,s292,s2721);
  and x331(s2750,s288,s2721);
  and x332(s2752,s280,s2721);
  and x333(s2754,s272,s2721);
  and x334(s2756,s264,s2721);
  and x335(s2758,s241,s2734);
  and x336(s2760,s233,s2734);
  and x337(s2762,s225,s2734);
  and x338(s2764,s217,s2734);
  and x339(s2766,s209,s2734);
  buf x340(s2827,s1701);
  not x341(s2838,s2828);
  not x342(s2847,s2822);
  not x343(s2885,s2882);
  not x344(s2889,s2886);
  not x345(s2893,s2890);
  not x346(s2897,s2894);
  not x347(s2901,s2898);
  not x348(s2905,s2902);
  and x349(s2906,s2393,s2886);
  and x350(s2909,s2393,s479,s2894);
  and x351(s2913,s2393,s490,s2902);
  and x352(s2918,s3554,s2882);
  and x353(s2922,s3554,s2890);
  and x354(s2927,s3554,s2898);
  not x355(s2951,s2948);
  not x356(s2955,s2952);
  not x357(s2959,s2956);
  not x358(s2963,s2960);
  not x359(s2967,s2964);
  not x360(s2971,s2968);
  and x361(s2973,s3553,s503,s2952);
  not x362(s2980,s2979);
  and x363(s2982,s3553,s523,s2960);
  and x364(s2988,s3553,s534,s2968);
  and x365(s2994,s3547,s2948);
  and x366(s3001,s3547,s2956);
  and x367(s3006,s3547,s2964);
  not x368(s3027,s3024);
  not x369(s3031,s3028);
  not x370(s3035,s3032);
  not x371(s3039,s3036);
  not x372(s3043,s3040);
  not x373(s3047,s3044);
  not x374(s3051,s3048);
  not x375(s3055,s3052);
  and x376(s3056,s2393,s389,s3028);
  and x377(s3060,s2393,s400,s3036);
  and x378(s3064,s2393,s411,s3044);
  and x379(s3068,s2393,s374,s3052);
  and x380(s3073,s3554,s3024);
  and x381(s3078,s3554,s3032);
  and x382(s3083,s3554,s3040);
  and x383(s3088,s3554,s3048);
  not x384(s3099,s3092);
  not x385(s3112,s3105);
  and x386(s3119,s372,s3092);
  and x387(s3121,s366,s3092);
  and x388(s3123,s358,s3092);
  and x389(s3125,s348,s3092);
  and x390(s3126,s338,s3092);
  and x391(s3128,s331,s3105);
  and x392(s3130,s323,s3105);
  and x393(s3132,s315,s3105);
  and x394(s3134,s307,s3105);
  and x395(s3136,s299,s3105);
  not x396(s3187,s3181);
  and x397(s3193,s83,s3181);
  and x398(s3196,s86,s3181);
  and x399(s3199,s88,s3181);
  and x400(s3202,s88,s3181);
  not x401(s3207,s3204);
  not x402(s3211,s3208);
  not x403(s3215,s3212);
  not x404(s3219,s3216);
  not x405(s3223,s3220);
  not x406(s3227,s3224);
  and x407(s3228,s2405,s503,s3208);
  and x408(s3232,s2405,s514);
  and x409(s3234,s2405,s523,s3216);
  and x410(s3238,s2405,s534,s3224);
  and x411(s3243,s3555,s3204);
  or x412(s3247,s3555,s514);
  and x413(s3249,s3555,s3212);
  and x414(s3253,s3555,s3220);
  not x415(s3259,s3256);
  not x416(s3263,s3260);
  not x417(s3267,s3264);
  not x418(s3271,s3268);
  not x419(s3275,s3272);
  not x420(s3279,s3276);
  and x421(s3280,s2405,s3260);
  and x422(s3283,s2405,s479,s3268);
  and x423(s3287,s2405,s490,s3276);
  and x424(s3292,s3555,s3256);
  and x425(s3295,s3555,s3264);
  and x426(s3299,s3555,s3272);
  not x427(s3305,s3302);
  buf x428(s3306,s2816);
  buf x429(s3310,s2816);
  not x430(s3317,s3314);
  buf x431(s3318,s2816);
  buf x432(s3322,s2816);
  and x433(s3326,s2405,s3302);
  and x434(s3333,s2405,s3314);
  not x435(s3357,s3354);
  not x436(s3361,s3358);
  not x437(s3365,s3362);
  not x438(s3369,s3366);
  not x439(s3373,s3370);
  not x440(s3377,s3374);
  not x441(s3381,s3378);
  not x442(s3385,s3382);
  and x443(s3386,s2393,s457,s3358);
  and x444(s3390,s2393,s468,s3366);
  and x445(s3394,s2393,s422,s3374);
  and x446(s3398,s2393,s435,s3382);
  and x447(s3403,s3554,s3354);
  and x448(s3408,s3554,s3362);
  and x449(s3413,s3554,s3370);
  and x450(s3418,s3554,s3378);
  not x451(s5088,s5082);
  not x452(s5089,s5085);
  not x453(s5096,s5090);
  not x454(s5097,s5093);
  buf x455(s3489,s3440);
  buf x456(s3493,s3440);
  not x457(s3570,s3558);
  not x458(s3594,s3582);
  not x459(s3622,s3616);
  not x460(s3632,s3628);
  and x461(s3637,s97,s3616);
  and x462(s3640,s94,s3616);
  and x463(s3643,s97,s3616);
  and x464(s3646,s94,s3616);
  not x465(s3672,s3660);
  not x466(s3696,s3684);
  not x467(s3745,s3737);
  not x468(s3765,s3757);
  not x469(s3803,s3795);
  not x470(s3823,s3815);
  not x471(s5338,s5332);
  not x472(s5339,s5335);
  not x473(s5346,s5340);
  not x474(s5347,s5343);
  not x475(s5354,s5348);
  not x476(s5355,s5351);
  not x477(s3979,s3972);
  not x478(s3998,s3991);
  not x479(s4037,s4030);
  not x480(s4056,s4049);
  buf x481(s4094,s4110);
  not x482(s5104,s5098);
  not x483(s5105,s5101);
  not x484(s5114,s5108);
  not x485(s5115,s5111);
  not x486(s5362,s5356);
  not x487(s5363,s5359);
  buf x488(s5366,s2816);
  not x489(s5373,s5369);
  buf x490(s993,s1688);
  buf x491(s978,s1688);
  buf x492(s949,s1688);
  buf x493(s939,s1688);
  and x494(s2568,s457,s3551,s2540);
  and x495(s2574,s468,s3551,s2548);
  and x496(s2580,s422,s3551,s2556);
  and x497(s2586,s435,s3551,s2564);
  and x498(s2592,s3549,s2536);
  and x499(s2597,s3549,s2544);
  and x500(s2602,s3549,s2552);
  and x501(s2607,s3549,s2560);
  and x502(s2662,s389,s3551,s2634);
  and x503(s2668,s400,s3551,s2642);
  and x504(s2674,s411,s3551,s2650);
  and x505(s2680,s374,s3551,s2658);
  and x506(s2686,s3549,s2630);
  and x507(s2691,s3549,s2638);
  and x508(s2696,s3549,s2646);
  and x509(s2701,s3549,s2654);
  and x510(s2907,s2370,s2889);
  and x511(s2910,s479,s2370,s2897);
  and x512(s2914,s490,s2370,s2905);
  and x513(s2920,s3556,s2885);
  and x514(s2924,s3556,s2893);
  and x515(s2929,s3556,s2901);
  and x516(s2975,s503,s3551,s2955);
  and x517(s2984,s523,s3551,s2963);
  and x518(s2990,s534,s3551,s2971);
  and x519(s2996,s3549,s2951);
  and x520(s3003,s3549,s2959);
  and x521(s3008,s3549,s2967);
  and x522(s3015,s2980,s2999);
  and x523(s3057,s389,s2370,s3031);
  and x524(s3061,s400,s2370,s3039);
  and x525(s3065,s411,s2370,s3047);
  and x526(s3069,s374,s2370,s3055);
  and x527(s3075,s3556,s3027);
  and x528(s3080,s3556,s3035);
  and x529(s3085,s3556,s3043);
  and x530(s3090,s3556,s3051);
  and x531(s3229,s503,s2382,s3211);
  not x532(s3233,s3232);
  and x533(s3235,s523,s2382,s3219);
  and x534(s3239,s534,s2382,s3227);
  and x535(s3244,s2361,s3207);
  and x536(s3250,s2361,s3215);
  and x537(s3254,s2361,s3223);
  and x538(s3281,s2382,s3263);
  and x539(s3284,s479,s2382,s3271);
  and x540(s3288,s490,s2382,s3279);
  and x541(s3293,s2361,s3259);
  and x542(s3296,s2361,s3267);
  and x543(s3300,s2361,s3275);
  and x544(s3327,s2382,s3305);
  and x545(s3334,s2382,s3317);
  and x546(s3387,s457,s2370,s3361);
  and x547(s3391,s468,s2370,s3369);
  and x548(s3395,s422,s2370,s3377);
  and x549(s3399,s435,s2370,s3385);
  and x550(s3405,s3556,s3357);
  and x551(s3410,s3556,s3365);
  and x552(s3415,s3556,s3373);
  and x553(s3420,s3556,s3381);
  nand x554(s3422,s5085,s5088);
  nand x555(s3423,s5082,s5089);
  nand x556(s3431,s5093,s5096);
  nand x557(s3432,s5090,s5097);
  nand x558(s3895,s5335,s5338);
  nand x559(s3896,s5332,s5339);
  nand x560(s3904,s5343,s5346);
  nand x561(s3905,s5340,s5347);
  nand x562(s3913,s5351,s5354);
  nand x563(s3914,s5348,s5355);
  buf x564(s889,s4094);
  nand x565(s5106,s5101,s5104);
  nand x566(s5107,s5098,s5105);
  nand x567(s5116,s5111,s5114);
  nand x568(s5117,s5108,s5115);
  nand x569(s5364,s5359,s5362);
  nand x570(s5365,s5356,s5363);
  not x571(s593,s4094);
  and x572(s2880,s2838,s2847);
  and x573(s2881,s2828,s2847);
  and x574(s1579,s200,s1540,s1552);
  and x575(s1585,s203,s1540,s1552);
  and x576(s1591,s197,s1540,s1552);
  and x577(s1597,s194,s1540,s1552);
  and x578(s1603,s191,s1540,s1552);
  and x579(s1667,s182,s1621,s1633);
  and x580(s1673,s188,s1621,s1633);
  and x581(s1679,s155,s1621,s1633);
  and x582(s1685,s149,s1621,s1633);
  and x583(s2876,s2838,s2847);
  and x584(s2877,s2828,s2847);
  and x585(s2253,s200,s2215,s2226);
  and x586(s2259,s203,s2215,s2226);
  and x587(s2265,s197,s2215,s2226);
  and x588(s2271,s194,s2215,s2226);
  and x589(s2277,s191,s2215,s2226);
  and x590(s2338,s182,s2293,s2304);
  and x591(s2344,s188,s2293,s2304);
  and x592(s2350,s155,s2293,s2304);
  and x593(s2356,s149,s2293,s2304);
  and x594(s2868,s2838,s2847);
  and x595(s2869,s2828,s2847);
  and x596(s710,s109,s3672,s3684);
  and x597(s2872,s2838,s2847);
  and x598(s2873,s2828,s2847);
  and x599(s720,s11,s2430,s2442);
  and x600(s725,s109,s3570,s3582);
  and x601(s730,s46,s3570,s3582);
  and x602(s735,s100,s3570,s3582);
  and x603(s740,s91,s3570,s3582);
  and x604(s745,s43,s3570,s3582);
  and x605(s750,s76,s2430,s2442);
  and x606(s755,s73,s2430,s2442);
  and x607(s760,s67,s2430,s2442);
  and x608(s765,s14,s2430,s2442);
  and x609(s770,s46,s3672,s3684);
  and x610(s775,s100,s3672,s3684);
  and x611(s780,s91,s3672,s3684);
  and x612(s785,s43,s3672,s3684);
  and x613(s790,s76,s2488,s2500);
  and x614(s795,s73,s2488,s2500);
  and x615(s800,s67,s2488,s2500);
  and x616(s805,s14,s2488,s2500);
  and x617(s841,s120,s3803,s3815);
  and x618(s857,s11,s2488,s2500);
  and x619(s880,s118,s3745,s3757);
  and x620(s1660,s176,s1621,s1633);
  and x621(s2331,s176,s2293,s2304);
  or x622(s2569,s2566,s2568);
  or x623(s2575,s2572,s2574);
  or x624(s2581,s2578,s2580);
  or x625(s2587,s2584,s2586);
  or x626(s2593,s2590,s2592,s457);
  or x627(s2598,s2595,s2597,s468);
  or x628(s2603,s2600,s2602,s422);
  or x629(s2608,s2605,s2607,s435);
  or x630(s2663,s2660,s2662);
  or x631(s2669,s2666,s2668);
  or x632(s2675,s2672,s2674);
  or x633(s2681,s2678,s2680);
  or x634(s2687,s2684,s2686,s389);
  or x635(s2692,s2689,s2691,s400);
  or x636(s2697,s2694,s2696,s411);
  or x637(s2702,s2699,s2701,s374);
  and x638(s2747,s289,s2728);
  and x639(s2749,s281,s2728);
  and x640(s2751,s273,s2728);
  and x641(s2753,s265,s2728);
  and x642(s2755,s257,s2728);
  and x643(s2757,s234,s2741);
  and x644(s2759,s226,s2741);
  and x645(s2761,s218,s2741);
  and x646(s2763,s210,s2741);
  and x647(s2765,s206,s2741);
  not x648(s2857,s2847);
  or x649(s2908,s2906,s2907);
  or x650(s2911,s2909,s2910);
  or x651(s2915,s2913,s2914);
  or x652(s2925,s2922,s2924,s479);
  or x653(s2930,s2927,s2929,s490);
  or x654(s2933,s2918,s2920);
  or x655(s2976,s2973,s2975);
  or x656(s2985,s2982,s2984);
  or x657(s2991,s2988,s2990);
  or x658(s2997,s2994,s2996,s503);
  or x659(s3004,s3001,s3003,s523);
  or x660(s3009,s3006,s3008,s534);
  or x661(s3058,s3056,s3057);
  or x662(s3062,s3060,s3061);
  or x663(s3066,s3064,s3065);
  or x664(s3070,s3068,s3069);
  or x665(s3076,s3073,s3075,s389);
  or x666(s3081,s3078,s3080,s400);
  or x667(s3086,s3083,s3085,s411);
  or x668(s3091,s3088,s3090,s374);
  and x669(s3118,s369,s3099);
  and x670(s3120,s361,s3099);
  and x671(s3122,s351,s3099);
  and x672(s3124,s341,s3099);
  and x673(s3127,s324,s3112);
  and x674(s3129,s316,s3112);
  and x675(s3131,s308,s3112);
  and x676(s3133,s302,s3112);
  and x677(s3135,s293,s3112);
  or x678(s3147,s3099,s3126);
  and x679(s3192,s83,s3187);
  and x680(s3195,s87,s3187);
  and x681(s3198,s34,s3187);
  and x682(s3201,s34,s3187);
  or x683(s3230,s3228,s3229);
  or x684(s3236,s3234,s3235);
  or x685(s3240,s3238,s3239);
  or x686(s3245,s3243,s3244,s503);
  or x687(s3251,s3249,s3250,s523);
  or x688(s3255,s3253,s3254,s534);
  or x689(s3282,s3280,s3281);
  or x690(s3285,s3283,s3284);
  or x691(s3289,s3287,s3288);
  or x692(s3297,s3295,s3296,s479);
  or x693(s3301,s3299,s3300,s490);
  not x694(s3309,s3306);
  not x695(s3313,s3310);
  not x696(s3321,s3318);
  not x697(s3325,s3322);
  or x698(s3328,s3326,s3327);
  and x699(s3329,s2405,s446,s3310);
  or x700(s3335,s3333,s3334);
  and x701(s3336,s2405,s446,s3322);
  and x702(s3341,s3555,s3306);
  and x703(s3345,s3555,s3318);
  or x704(s3388,s3386,s3387);
  or x705(s3392,s3390,s3391);
  or x706(s3396,s3394,s3395);
  or x707(s3400,s3398,s3399);
  or x708(s3406,s3403,s3405,s457);
  or x709(s3411,s3408,s3410,s468);
  or x710(s3416,s3413,s3415,s422);
  or x711(s3421,s3418,s3420,s435);
  nand x712(s3424,s3422,s3423);
  nand x713(s3433,s3431,s3432);
  not x714(s3492,s3489);
  not x715(s3496,s3493);
  and x716(s3780,s117,s3745,s3757);
  and x717(s3783,s126,s3745,s3757);
  and x718(s3786,s127,s3745,s3757);
  and x719(s3789,s128,s3745,s3757);
  and x720(s3838,s131,s3803,s3815);
  and x721(s3841,s129,s3803,s3815);
  and x722(s3844,s119,s3803,s3815);
  and x723(s3847,s130,s3803,s3815);
  nand x724(s3897,s3895,s3896);
  nand x725(s3906,s3904,s3905);
  nand x726(s3915,s3913,s3914);
  and x727(s4011,s122,s3979,s3991);
  and x728(s4014,s113,s3979,s3991);
  and x729(s4017,s53,s3979,s3991);
  and x730(s4020,s114,s3979,s3991);
  and x731(s4023,s115,s3979,s3991);
  and x732(s4069,s52,s4037,s4049);
  and x733(s4072,s112,s4037,s4049);
  and x734(s4075,s116,s4037,s4049);
  and x735(s4078,s121,s4037,s4049);
  and x736(s4081,s123,s4037,s4049);
  nand x737(s5206,s5116,s5117);
  nand x738(s5209,s5106,s5107);
  and x739(s5307,s3233,s3247);
  or x740(s5322,s3292,s3293);
  not x741(s5372,s5366);
  nand x742(s5375,s5366,s5373);
  nand x743(s5399,s5364,s5365);
  not x744(s2813,s3015);
  or x745(s3197,s3195,s3196);
  or x746(s3200,s3198,s3199);
  or x747(s3203,s3201,s3202);
  or x748(s3194,s3192,s3193);
  not x749(s2570,s2569);
  not x750(s2576,s2575);
  not x751(s2582,s2581);
  not x752(s2588,s2587);
  not x753(s2664,s2663);
  not x754(s2670,s2669);
  not x755(s2676,s2675);
  not x756(s2682,s2681);
  or x757(s2767,s2749,s2750);
  or x758(s2772,s2751,s2752);
  or x759(s2776,s2753,s2754);
  or x760(s2780,s2755,s2756);
  or x761(s2784,s2757,s2758);
  or x762(s2788,s2759,s2760);
  or x763(s2794,s2761,s2762);
  or x764(s2798,s2763,s2764);
  or x765(s2802,s2765,s2766);
  not x766(s2912,s2911);
  not x767(s2916,s2915);
  not x768(s2936,s2908);
  not x769(s2977,s2976);
  not x770(s2986,s2985);
  not x771(s2992,s2991);
  not x772(s3059,s3058);
  not x773(s3063,s3062);
  not x774(s3067,s3066);
  not x775(s3071,s3070);
  or x776(s3137,s3120,s3121);
  or x777(s3139,s3122,s3123);
  or x778(s3143,s3124,s3125);
  or x779(s3151,s3127,s3128);
  or x780(s3155,s3129,s3130);
  or x781(s3161,s3131,s3132);
  or x782(s3165,s3133,s3134);
  or x783(s3167,s3135,s3136);
  not x784(s3231,s3230);
  not x785(s3237,s3236);
  not x786(s3241,s3240);
  not x787(s3286,s3285);
  not x788(s3290,s3289);
  and x789(s3330,s446,s2382,s3313);
  and x790(s3337,s446,s2382,s3325);
  and x791(s3342,s2361,s3309);
  and x792(s3346,s2361,s3321);
  not x793(s3348,s3328);
  not x794(s3352,s3335);
  not x795(s3389,s3388);
  not x796(s3393,s3392);
  not x797(s3397,s3396);
  not x798(s3401,s3400);
  and x799(s3845,s3015,s3803,s3823);
  or x800(s5126,s3118,s3119);
  or x801(s5178,s2747,s2748);
  not x802(s5325,s3282);
  nand x803(s5374,s5369,s5372);
  not x804(s2810,s2933);
  and x805(s635,s3197,s3176);
  and x806(s2878,s24,s2838,s2857);
  and x807(s2879,s25,s2828,s2857);
  and x808(s2874,s26,s2838,s2857);
  and x809(s2875,s81,s2828,s2857);
  and x810(s703,s3200,s3176);
  and x811(s2866,s79,s2838,s2857);
  and x812(s2867,s23,s2828,s2857);
  and x813(s2870,s82,s2838,s2857);
  and x814(s2871,s80,s2828,s2857);
  and x815(s716,s3203,s3176);
  and x816(s819,s3194,s3176);
  and x817(s1789,s3147,s514);
  and x818(s2036,s514,s3147);
  and x819(s2611,s2570,s2593);
  and x820(s2615,s2576,s2598);
  and x821(s2619,s2582,s2603);
  and x822(s2623,s2588,s2608);
  and x823(s2705,s2664,s2687);
  and x824(s2709,s2670,s2692);
  and x825(s2713,s2676,s2697);
  and x826(s2717,s2682,s2702);
  and x827(s2939,s2912,s2925);
  and x828(s2942,s2916,s2930);
  buf x829(s2945,s2933);
  and x830(s3012,s2977,s2997);
  and x831(s3018,s2986,s3004);
  and x832(s3021,s2992,s3009);
  or x833(s3331,s3329,s3330);
  or x834(s3338,s3336,s3337);
  or x835(s3343,s3341,s3342,s446);
  or x836(s3347,s3345,s3346,s446);
  not x837(s3428,s3424);
  not x838(s3437,s3433);
  and x839(s3514,s3433,s3424,s3489);
  and x840(s3836,s3352,s3803,s3823);
  and x841(s3852,s3071,s3091);
  not x842(s5311,s5307);
  not x843(s3901,s3897);
  not x844(s3910,s3906);
  buf x845(s3934,s3915);
  buf x846(s3938,s3915);
  buf x847(s4652,s3147);
  buf x848(s4783,s3147);
  buf x849(s5137,s3147);
  not x850(s5212,s5206);
  not x851(s5213,s5209);
  and x852(s5260,s3063,s3081);
  and x853(s5263,s3067,s3086);
  and x854(s5268,s3401,s3421);
  and x855(s5271,s3059,s3076);
  and x856(s5276,s3393,s3411);
  and x857(s5279,s3397,s3416);
  and x858(s5289,s3389,s3406);
  and x859(s5296,s3237,s3251);
  and x860(s5299,s3241,s3255);
  and x861(s5304,s3231,s3245);
  and x862(s5312,s3286,s3297);
  and x863(s5315,s3290,s3301);
  not x864(s5328,s5322);
  nand x865(s5396,s5374,s5375);
  not x866(s5403,s5399);
  and x867(s1286,s446,s2802);
  not x868(s2809,s2936);
  not x869(s597,s3348);
  and x870(s1031,s2802,s446);
  not x871(s636,s635);
  or x872(s637,s2878,s2879,s2880,s2881);
  or x873(s671,s2874,s2875,s2876,s2877);
  not x874(s704,s703);
  or x875(s705,s2866,s2867,s2868,s2869);
  or x876(s713,s2870,s2871,s2872,s2873);
  not x877(s717,s716);
  not x878(s820,s819);
  and x879(s1046,s2798,s457);
  and x880(s1064,s2794,s468);
  and x881(s1071,s422,s2788);
  and x882(s1097,s2784,s435);
  and x883(s1111,s2780,s389);
  and x884(s1128,s2776,s400);
  and x885(s1145,s2772,s411);
  and x886(s1160,s2767,s374);
  and x887(s1301,s457,s2798);
  and x888(s1318,s468,s2794);
  and x889(s1324,s422,s2788);
  and x890(s1341,s435,s2784);
  and x891(s1359,s389,s2780);
  and x892(s1382,s400,s2776);
  and x893(s1404,s411,s2772);
  and x894(s1412,s374,s2767);
  not x895(s1704,s3167);
  not x896(s1712,s3165);
  buf x897(s1724,s3165);
  and x898(s1742,s3161,s479);
  and x899(s1749,s490,s3155);
  and x900(s1775,s3151,s503);
  and x901(s1806,s3143,s523);
  and x902(s1823,s3139,s534);
  not x903(s1829,s3137);
  buf x904(s1837,s3137);
  not x905(s1958,s3167);
  not x906(s1966,s3165);
  buf x907(s1978,s3165);
  and x908(s1995,s479,s3161);
  and x909(s2001,s490,s3155);
  and x910(s2018,s503,s3151);
  and x911(s2059,s523,s3143);
  and x912(s2081,s534,s3139);
  buf x913(s2089,s3137);
  not x914(s2106,s3137);
  buf x915(s3170,s3167);
  not x916(s3332,s3331);
  not x917(s3339,s3338);
  not x918(s5132,s5126);
  not x919(s5184,s5178);
  not x920(s3853,s3852);
  not x921(s3874,s3348);
  and x922(s4076,s2936,s4037,s4056);
  buf x923(s4116,s2802);
  buf x924(s4124,s2798);
  buf x925(s4132,s2794);
  buf x926(s4140,s2788);
  buf x927(s4148,s2784);
  buf x928(s4156,s2780);
  buf x929(s4164,s2776);
  buf x930(s4172,s2772);
  buf x931(s4180,s2767);
  nor x932(s4228,s422,s2788);
  buf x933(s4279,s2802);
  buf x934(s4287,s2798);
  buf x935(s4295,s2794);
  buf x936(s4303,s2784);
  buf x937(s4311,s2780);
  buf x938(s4319,s2776);
  buf x939(s4327,s2772);
  buf x940(s4335,s2788);
  buf x941(s4343,s2767);
  nor x942(s4348,s422,s2788);
  nor x943(s4464,s374,s2767);
  buf x944(s4628,s3161);
  buf x945(s4636,s3155);
  buf x946(s4644,s3151);
  buf x947(s4660,s3143);
  buf x948(s4668,s3139);
  nor x949(s4716,s490,s3155);
  buf x950(s4767,s3161);
  buf x951(s4775,s3151);
  buf x952(s4791,s3143);
  buf x953(s4799,s3139);
  buf x954(s4807,s3155);
  nor x955(s4812,s490,s3155);
  buf x956(s5118,s3139);
  buf x957(s5121,s3143);
  buf x958(s5129,s3137);
  buf x959(s5134,s3151);
  buf x960(s5142,s3161);
  buf x961(s5145,s3155);
  buf x962(s5152,s3167);
  buf x963(s5155,s3165);
  buf x964(s5162,s2788);
  buf x965(s5165,s2784);
  buf x966(s5170,s2798);
  buf x967(s5173,s2794);
  buf x968(s5181,s2802);
  buf x969(s5186,s2772);
  buf x970(s5189,s2767);
  buf x971(s5196,s2780);
  buf x972(s5199,s2776);
  nand x973(s5214,s5209,s5212);
  nand x974(s5215,s5206,s5213);
  not x975(s5329,s5325);
  nand x976(s5330,s5325,s5328);
  not x977(s2807,s2942);
  not x978(s2808,s2939);
  not x979(s2811,s3021);
  not x980(s2812,s3018);
  not x981(s2814,s3012);
  not x982(s2626,s2623);
  not x983(s2622,s2619);
  not x984(s2618,s2615);
  not x985(s2614,s2611);
  not x986(s2720,s2717);
  not x987(s2716,s2713);
  not x988(s2712,s2709);
  not x989(s2708,s2705);
  and x990(s639,s637,s2827);
  and x991(s673,s671,s2827);
  and x992(s707,s705,s2827);
  and x993(s715,s713,s2827);
  and x994(s3731,s2945,s3728,s3721);
  not x995(s4658,s4652);
  nand x996(s1777,s4652,s4659);
  nand x997(s2019,s4783,s4786);
  not x998(s4787,s4783);
  and x999(s3350,s3332,s3343);
  and x1000(s3353,s3339,s3347);
  not x1001(s5141,s5137);
  and x1002(s3513,s3428,s3433,s3492);
  and x1003(s3516,s3424,s3437,s3496);
  and x1004(s3517,s3437,s3428,s3493);
  and x1005(s3778,s2717,s3745,s3765);
  and x1006(s3781,s2713,s3745,s3765);
  and x1007(s3784,s2709,s3745,s3765);
  and x1008(s3787,s2705,s3745,s3765);
  and x1009(s3839,s3021,s3803,s3823);
  and x1010(s3842,s3018,s3803,s3823);
  not x1011(s5266,s5260);
  not x1012(s5267,s5263);
  not x1013(s5274,s5268);
  not x1014(s5275,s5271);
  not x1015(s5302,s5296);
  not x1016(s5303,s5299);
  not x1017(s5310,s5304);
  nand x1018(s3891,s5304,s5311);
  not x1019(s3937,s3934);
  not x1020(s3941,s3938);
  and x1021(s3955,s3906,s3897,s3934);
  and x1022(s3958,s3910,s3901,s3938);
  and x1023(s4009,s2623,s3979,s3998);
  and x1024(s4012,s2619,s3979,s3998);
  and x1025(s4015,s2615,s3979,s3998);
  and x1026(s4018,s2611,s3979,s3998);
  and x1027(s4067,s3012,s4037,s4056);
  and x1028(s4070,s2942,s4037,s4056);
  and x1029(s4073,s2939,s4037,s4056);
  and x1030(s4079,s2945,s4037,s4056);
  nand x1031(s5239,s5214,s5215);
  not x1032(s5282,s5276);
  not x1033(s5283,s5279);
  not x1034(s5293,s5289);
  not x1035(s5318,s5312);
  not x1036(s5319,s5315);
  nand x1037(s5331,s5322,s5329);
  not x1038(s5402,s5396);
  nand x1039(s5405,s5396,s5403);
  and x1040(s595,s2807,s2808,s2809,s2810);
  and x1041(s596,s2811,s2812,s2813,s2814);
  and x1042(s607,s2626,s2622,s2618,s2614);
  and x1043(s608,s2720,s2716,s2712,s2708);
  and x1044(s1845,s1704,s1724);
  and x1045(s1846,s1712,s1704,s1742);
  and x1046(s2115,s1958,s1978);
  and x1047(s2116,s1966,s1958,s1995);
  not x1048(s4122,s4116);
  nand x1049(s1022,s4116,s4123);
  not x1050(s4130,s4124);
  nand x1051(s1033,s4124,s4131);
  not x1052(s4138,s4132);
  nand x1053(s1051,s4132,s4139);
  not x1054(s4146,s4140);
  nand x1055(s1079,s4140,s4147);
  not x1056(s4154,s4148);
  nand x1057(s1088,s4148,s4155);
  not x1058(s4162,s4156);
  nand x1059(s1099,s4156,s4163);
  not x1060(s4170,s4164);
  nand x1061(s1115,s4164,s4171);
  not x1062(s4178,s4172);
  nand x1063(s1133,s4172,s4179);
  not x1064(s4186,s4180);
  nand x1065(s1151,s4180,s4187);
  not x1066(s4234,s4228);
  nand x1067(s1276,s4279,s4282);
  not x1068(s4283,s4279);
  nand x1069(s1287,s4287,s4290);
  not x1070(s4291,s4287);
  nand x1071(s1305,s4295,s4298);
  not x1072(s4299,s4295);
  nand x1073(s1330,s4303,s4306);
  not x1074(s4307,s4303);
  nand x1075(s1342,s4311,s4314);
  not x1076(s4315,s4311);
  nand x1077(s1363,s4319,s4322);
  not x1078(s4323,s4319);
  nand x1079(s1388,s4327,s4330);
  not x1080(s4331,s4327);
  nand x1081(s1420,s4335,s4338);
  not x1082(s4339,s4335);
  nand x1083(s1428,s4343,s4346);
  not x1084(s4347,s4343);
  not x1085(s4634,s4628);
  nand x1086(s1729,s4628,s4635);
  not x1087(s4642,s4636);
  nand x1088(s1757,s4636,s4643);
  not x1089(s4650,s4644);
  nand x1090(s1766,s4644,s4651);
  nand x1091(s1776,s4655,s4658);
  not x1092(s4666,s4660);
  nand x1093(s1793,s4660,s4667);
  not x1094(s4674,s4668);
  nand x1095(s1811,s4668,s4675);
  and x1096(s1849,s1712,s1742);
  and x1097(s1852,s1712,s1742);
  and x1098(s1875,s54,s1829);
  not x1099(s4722,s4716);
  nand x1100(s1982,s4767,s4770);
  not x1101(s4771,s4767);
  nand x1102(s2007,s4775,s4778);
  not x1103(s4779,s4775);
  nand x1104(s2020,s4780,s4787);
  nand x1105(s2040,s4791,s4794);
  not x1106(s4795,s4791);
  nand x1107(s2065,s4799,s4802);
  not x1108(s4803,s4799);
  nand x1109(s2097,s4807,s4810);
  not x1110(s4811,s4807);
  and x1111(s2119,s1966,s1995);
  and x1112(s2122,s1966,s1995);
  not x1113(s5124,s5118);
  not x1114(s5125,s5121);
  nand x1115(s3452,s5129,s5132);
  not x1116(s5133,s5129);
  not x1117(s5140,s5134);
  nand x1118(s3462,s5134,s5141);
  not x1119(s5168,s5162);
  not x1120(s5169,s5165);
  not x1121(s5176,s5170);
  not x1122(s5177,s5173);
  nand x1123(s3484,s5181,s5184);
  not x1124(s5185,s5181);
  nor x1125(s3515,s3513,s3514);
  nor x1126(s3518,s3516,s3517);
  not x1127(s3857,s3853);
  nand x1128(s3860,s5263,s5266);
  nand x1129(s3861,s5260,s5267);
  nand x1130(s3869,s5271,s5274);
  nand x1131(s3870,s5268,s5275);
  not x1132(s3878,s3874);
  nand x1133(s3881,s5299,s5302);
  nand x1134(s3882,s5296,s5303);
  nand x1135(s3890,s5307,s5310);
  and x1136(s3954,s3901,s3906,s3937);
  and x1137(s3957,s3897,s3910,s3941);
  and x1138(s4021,s3353,s3979,s3998);
  not x1139(s4099,s3170);
  buf x1140(s4236,s1071);
  not x1141(s4354,s4348);
  buf x1142(s4406,s1324);
  not x1143(s4470,s4464);
  buf x1144(s4552,s1412);
  buf x1145(s4679,s1829);
  buf x1146(s4687,s1704);
  buf x1147(s4695,s1704);
  buf x1148(s4703,s1712);
  buf x1149(s4711,s1712);
  buf x1150(s4724,s1749);
  not x1151(s4818,s4812);
  buf x1152(s4855,s1958);
  buf x1153(s4865,s1966);
  buf x1154(s4870,s2001);
  buf x1155(s4913,s1958);
  buf x1156(s4923,s1966);
  buf x1157(s4951,s2106);
  buf x1158(s5006,s2089);
  buf x1159(s5039,s2106);
  not x1160(s5148,s5142);
  not x1161(s5149,s5145);
  not x1162(s5158,s5152);
  not x1163(s5159,s5155);
  not x1164(s5192,s5186);
  not x1165(s5193,s5189);
  not x1166(s5202,s5196);
  not x1167(s5203,s5199);
  nand x1168(s5284,s5279,s5282);
  nand x1169(s5285,s5276,s5283);
  nand x1170(s5320,s5315,s5318);
  nand x1171(s5321,s5312,s5319);
  nand x1172(s5386,s5330,s5331);
  nand x1173(s5404,s5399,s5402);
  and x1174(s598,s595,s596,s597);
  not x1175(s609,s3350);
  nand x1176(s1021,s4119,s4122);
  nand x1177(s1032,s4127,s4130);
  nand x1178(s1050,s4135,s4138);
  nand x1179(s1078,s4143,s4146);
  nand x1180(s1087,s4151,s4154);
  nand x1181(s1098,s4159,s4162);
  nand x1182(s1114,s4167,s4170);
  nand x1183(s1132,s4175,s4178);
  nand x1184(s1150,s4183,s4186);
  nand x1185(s1277,s4276,s4283);
  nand x1186(s1288,s4284,s4291);
  nand x1187(s1306,s4292,s4299);
  nand x1188(s1331,s4300,s4307);
  nand x1189(s1343,s4308,s4315);
  nand x1190(s1364,s4316,s4323);
  nand x1191(s1389,s4324,s4331);
  nand x1192(s1421,s4332,s4339);
  nand x1193(s1429,s4340,s4347);
  nand x1194(s1728,s4631,s4634);
  nand x1195(s1756,s4639,s4642);
  nand x1196(s1765,s4647,s4650);
  nand x1197(s1778,s1776,s1777);
  nand x1198(s1792,s4663,s4666);
  nand x1199(s1810,s4671,s4674);
  nand x1200(s1983,s4764,s4771);
  nand x1201(s2008,s4772,s4779);
  nand x1202(s2021,s2019,s2020);
  nand x1203(s2041,s4788,s4795);
  nand x1204(s2066,s4796,s4803);
  nand x1205(s2098,s4804,s4811);
  nand x1206(s3443,s5121,s5124);
  nand x1207(s3444,s5118,s5125);
  nand x1208(s3453,s5126,s5133);
  nand x1209(s3461,s5137,s5140);
  nand x1210(s3466,s5165,s5168);
  nand x1211(s3467,s5162,s5169);
  nand x1212(s3475,s5173,s5176);
  nand x1213(s3476,s5170,s5177);
  nand x1214(s3485,s5178,s5185);
  not x1215(s5243,s5239);
  nand x1216(s3862,s3860,s3861);
  nand x1217(s3871,s3869,s3870);
  nand x1218(s3883,s3881,s3882);
  nand x1219(s3892,s3890,s3891);
  nor x1220(s3956,s3954,s3955);
  nor x1221(s3959,s3957,s3958);
  or x1222(s4756,s1837,s1875);
  nand x1223(s5150,s5145,s5148);
  nand x1224(s5151,s5142,s5149);
  nand x1225(s5160,s5155,s5158);
  nand x1226(s5161,s5152,s5159);
  nand x1227(s5194,s5189,s5192);
  nand x1228(s5195,s5186,s5193);
  nand x1229(s5204,s5199,s5202);
  nand x1230(s5205,s5196,s5203);
  nand x1231(s5236,s3518,s3515);
  buf x1232(s5286,s3350);
  nand x1233(s5379,s5284,s5285);
  nand x1234(s5389,s5320,s5321);
  nand x1235(s5425,s5404,s5405);
  and x1236(s610,s607,s608,s609);
  nand x1237(s1023,s1021,s1022);
  nand x1238(s1034,s1032,s1033);
  nand x1239(s1052,s1050,s1051);
  nand x1240(s1080,s1078,s1079);
  nand x1241(s1089,s1087,s1088);
  nand x1242(s1100,s1098,s1099);
  nand x1243(s1116,s1114,s1115);
  nand x1244(s1134,s1132,s1133);
  nand x1245(s1152,s1150,s1151);
  not x1246(s4242,s4236);
  nand x1247(s1278,s1276,s1277);
  nand x1248(s1289,s1287,s1288);
  nand x1249(s1307,s1305,s1306);
  nand x1250(s1332,s1330,s1331);
  nand x1251(s1344,s1342,s1343);
  nand x1252(s1365,s1363,s1364);
  nand x1253(s1390,s1388,s1389);
  nand x1254(s1422,s1420,s1421);
  nand x1255(s1430,s1428,s1429);
  nand x1256(s1730,s1728,s1729);
  nand x1257(s1758,s1756,s1757);
  nand x1258(s1767,s1765,s1766);
  nand x1259(s1794,s1792,s1793);
  nand x1260(s1812,s1810,s1811);
  nand x1261(s1876,s4679,s4682);
  not x1262(s4683,s4679);
  not x1263(s4691,s4687);
  not x1264(s4699,s4695);
  not x1265(s4707,s4703);
  not x1266(s4715,s4711);
  not x1267(s4730,s4724);
  nand x1268(s1984,s1982,s1983);
  nand x1269(s2009,s2007,s2008);
  nand x1270(s2042,s2040,s2041);
  nand x1271(s2067,s2065,s2066);
  nand x1272(s2099,s2097,s2098);
  not x1273(s4869,s4865);
  not x1274(s4927,s4923);
  nand x1275(s3445,s3443,s3444);
  nand x1276(s3454,s3452,s3453);
  nand x1277(s3463,s3461,s3462);
  nand x1278(s3468,s3466,s3467);
  nand x1279(s3477,s3475,s3476);
  nand x1280(s3486,s3484,s3485);
  and x1281(s4103,s4099,s3170);
  not x1282(s4412,s4406);
  not x1283(s4558,s4552);
  not x1284(s4859,s4855);
  not x1285(s4876,s4870);
  not x1286(s4917,s4913);
  not x1287(s4955,s4951);
  not x1288(s5012,s5006);
  not x1289(s5043,s5039);
  nand x1290(s5216,s5160,s5161);
  nand x1291(s5219,s5150,s5151);
  nand x1292(s5226,s5204,s5205);
  nand x1293(s5229,s5194,s5195);
  not x1294(s5392,s5386);
  nand x1295(s5422,s3959,s3956);
  and x1296(s1866,s1778,s1806);
  nand x1297(s1877,s4676,s4683);
  not x1298(s4762,s4756);
  and x1299(s2142,s2021,s2059);
  and x1300(s2146,s2021,s2059);
  not x1301(s5242,s5236);
  nand x1302(s3532,s5236,s5243);
  not x1303(s3866,s3862);
  not x1304(s3887,s3883);
  buf x1305(s3918,s3871);
  buf x1306(s3922,s3871);
  buf x1307(s3926,s3892);
  buf x1308(s3930,s3892);
  not x1309(s5429,s5425);
  or x1310(s4104,s4099,s4103);
  buf x1311(s4743,s1778);
  buf x1312(s4991,s2021);
  buf x1313(s5001,s2021);
  not x1314(s5292,s5286);
  nand x1315(s5295,s5286,s5293);
  not x1316(s5383,s5379);
  not x1317(s5393,s5389);
  nand x1318(s5394,s5389,s5392);
  and x1319(s1439,s1278,s1301);
  and x1320(s1440,s1289,s1278,s1318);
  and x1321(s1441,s1307,s1278,s1324,s1289);
  and x1322(s1847,s1730,s1704,s1749,s1712);
  and x1323(s1168,s1023,s1046);
  and x1324(s1169,s1034,s1023,s1064);
  and x1325(s1170,s1052,s1023,s1071,s1034);
  and x1326(s2117,s1984,s1958,s2001,s1966);
  not x1327(s1086,s1080);
  and x1328(s1166,s1034,s1080,s1052,s1023);
  and x1329(s1171,s1034,s1064);
  and x1330(s1172,s1052,s1071,s1034);
  and x1331(s1173,s1080,s1052,s1034);
  and x1332(s1174,s1034,s1064);
  and x1333(s1175,s1071,s1052,s1034);
  and x1334(s1176,s1052,s1071);
  and x1335(s1177,s1080,s1052);
  and x1336(s1178,s1052,s1071);
  and x1337(s1179,s1100,s1152,s1116,s1089,s1134);
  and x1338(s1181,s1089,s1111);
  and x1339(s1182,s1100,s1089,s1128);
  and x1340(s1183,s1116,s1089,s1145,s1100);
  and x1341(s1184,s1134,s1116,s1089,s1160,s1100);
  and x1342(s1188,s1100,s1128);
  and x1343(s1189,s1116,s1145,s1100);
  and x1344(s1190,s1134,s1116,s1160,s1100);
  and x1345(s1191,s4,s1152,s1116,s1134,s1100);
  and x1346(s1192,s1145,s1116);
  and x1347(s1193,s1134,s1116,s1160);
  and x1348(s1194,s4,s1152,s1116,s1134);
  and x1349(s1195,s1134,s1160);
  and x1350(s1196,s4,s1152,s1134);
  and x1351(s1197,s4,s1152);
  and x1352(s1437,s1422,s1307,s1289,s1278);
  and x1353(s1442,s1289,s1318);
  and x1354(s1443,s1307,s1324,s1289);
  and x1355(s1444,s1422,s1307,s1289);
  and x1356(s1445,s1289,s1318);
  and x1357(s1446,s1307,s1324,s1289);
  and x1358(s1447,s1307,s1324);
  and x1359(s1451,s1430,s1390,s1365,s1344,s1332);
  and x1360(s1454,s1332,s1359);
  and x1361(s1455,s1344,s1332,s1382);
  and x1362(s1456,s1365,s1332,s1404,s1344);
  and x1363(s1457,s1390,s1365,s1332,s1412,s1344);
  and x1364(s1465,s1344,s1382);
  and x1365(s1466,s1365,s1404,s1344);
  and x1366(s1467,s1390,s1365,s1412,s1344);
  and x1367(s1468,s1430,s1365,s1344,s1390);
  and x1368(s1469,s1344,s1382);
  and x1369(s1470,s1365,s1404,s1344);
  and x1370(s1471,s1390,s1365,s1412,s1344);
  and x1371(s1472,s1365,s1404);
  and x1372(s1473,s1390,s1365,s1412);
  and x1373(s1474,s1430,s1365,s1390);
  and x1374(s1475,s1365,s1404);
  and x1375(s1476,s1390,s1365,s1412);
  and x1376(s1477,s1390,s1412);
  and x1377(s1481,s1422,s1307);
  and x1378(s1482,s1430,s1390);
  not x1379(s1764,s1758);
  and x1380(s1843,s1712,s1758,s1730,s1704);
  and x1381(s1850,s1730,s1749,s1712);
  and x1382(s1851,s1758,s1730,s1712);
  and x1383(s1853,s1749,s1730,s1712);
  and x1384(s1854,s1730,s1749);
  and x1385(s1855,s1758,s1730);
  and x1386(s1856,s1730,s1749);
  and x1387(s1857,s1778,s1829,s1794,s1767,s1812);
  and x1388(s1859,s1767,s1789);
  and x1389(s1860,s1778,s1767,s1806);
  and x1390(s1861,s1794,s1767,s1823,s1778);
  and x1391(s1862,s1812,s1794,s1767,s1837,s1778);
  and x1392(s1867,s1794,s1823,s1778);
  and x1393(s1868,s1812,s1794,s1837,s1778);
  and x1394(s1869,s54,s1829,s1794,s1812,s1778);
  and x1395(s1870,s1823,s1794);
  and x1396(s1871,s1812,s1794,s1837);
  and x1397(s1872,s54,s1829,s1794,s1812);
  and x1398(s1873,s1812,s1837);
  and x1399(s1874,s54,s1829,s1812);
  nand x1400(s1878,s1876,s1877);
  and x1401(s2113,s2099,s1984,s1966,s1958);
  and x1402(s2120,s1984,s2001,s1966);
  and x1403(s2121,s2099,s1984,s1966);
  and x1404(s2123,s1984,s2001,s1966);
  and x1405(s2124,s1984,s2001);
  and x1406(s2128,s2106,s2067,s2042,s2021,s2009);
  and x1407(s2131,s2009,s2036);
  and x1408(s2132,s2021,s2009,s2059);
  and x1409(s2133,s2042,s2009,s2081,s2021);
  and x1410(s2134,s2067,s2042,s2009,s2089,s2021);
  and x1411(s2143,s2042,s2081,s2021);
  and x1412(s2144,s2067,s2042,s2089,s2021);
  and x1413(s2145,s2106,s2042,s2021,s2067);
  and x1414(s2147,s2042,s2081,s2021);
  and x1415(s2148,s2067,s2042,s2089,s2021);
  and x1416(s2149,s2042,s2081);
  and x1417(s2150,s2067,s2042,s2089);
  and x1418(s2151,s2106,s2042,s2067);
  and x1419(s2152,s2042,s2081);
  and x1420(s2153,s2067,s2042,s2089);
  and x1421(s2154,s2067,s2089);
  and x1422(s2158,s2099,s1984);
  and x1423(s2159,s2106,s2067);
  not x1424(s3449,s3445);
  not x1425(s3458,s3454);
  not x1426(s3472,s3468);
  not x1427(s3481,s3477);
  buf x1428(s3497,s3463);
  buf x1429(s3501,s3463);
  buf x1430(s3505,s3486);
  buf x1431(s3509,s3486);
  nand x1432(s3531,s5239,s5242);
  not x1433(s5428,s5422);
  nand x1434(s3967,s5422,s5429);
  buf x1435(s4191,s1152);
  buf x1436(s4199,s1023);
  buf x1437(s4207,s1023);
  buf x1438(s4215,s1034);
  buf x1439(s4223,s1034);
  buf x1440(s4231,s1052);
  buf x1441(s4239,s1052);
  buf x1442(s4247,s1089);
  buf x1443(s4255,s1100);
  buf x1444(s4263,s1116);
  buf x1445(s4271,s1134);
  buf x1446(s4371,s1422);
  buf x1447(s4381,s1307);
  buf x1448(s4391,s1278);
  buf x1449(s4401,s1289);
  buf x1450(s4429,s1422);
  buf x1451(s4439,s1307);
  buf x1452(s4449,s1278);
  buf x1453(s4459,s1289);
  buf x1454(s4497,s1430);
  buf x1455(s4507,s1390);
  buf x1456(s4517,s1332);
  buf x1457(s4527,s1365);
  buf x1458(s4537,s1344);
  buf x1459(s4547,s1344);
  buf x1460(s4585,s1430);
  buf x1461(s4595,s1390);
  buf x1462(s4605,s1332);
  buf x1463(s4615,s1365);
  buf x1464(s4719,s1730);
  buf x1465(s4727,s1730);
  buf x1466(s4735,s1767);
  buf x1467(s4751,s1794);
  buf x1468(s4759,s1812);
  buf x1469(s4835,s2099);
  buf x1470(s4845,s1984);
  buf x1471(s4893,s2099);
  buf x1472(s4903,s1984);
  buf x1473(s4961,s2067);
  buf x1474(s4971,s2009);
  buf x1475(s4981,s2042);
  buf x1476(s5049,s2067);
  buf x1477(s5059,s2009);
  buf x1478(s5069,s2042);
  not x1479(s5222,s5216);
  not x1480(s5223,s5219);
  not x1481(s5232,s5226);
  not x1482(s5233,s5229);
  nand x1483(s5294,s5289,s5292);
  nand x1484(s5395,s5386,s5393);
  or x1485(s589,s1286,s1439,s1440,s1441);
  or x1486(s616,s3167,s1845,s1846,s1847);
  or x1487(s619,s1031,s1168,s1169,s1170);
  or x1488(s627,s3167,s2115,s2116,s2117);
  or x1489(s1185,s1097,s1181,s1182,s1183,s1184);
  or x1490(s1448,s1318,s1447);
  or x1491(s1458,s1341,s1454,s1455,s1456,s1457);
  or x1492(s1478,s1404,s1477);
  or x1493(s1863,s1775,s1859,s1860,s1861,s1862);
  not x1494(s4747,s4743);
  or x1495(s2125,s1995,s2124);
  or x1496(s2135,s2018,s2131,s2132,s2133,s2134);
  or x1497(s2155,s2081,s2154);
  not x1498(s4995,s4991);
  not x1499(s5005,s5001);
  nand x1500(s3533,s3531,s3532);
  not x1501(s3921,s3918);
  not x1502(s3925,s3922);
  not x1503(s3929,s3926);
  not x1504(s3933,s3930);
  and x1505(s3943,s3862,s3853,s3918);
  and x1506(s3946,s3866,s3857,s3922);
  and x1507(s3949,s3883,s3874,s3926);
  and x1508(s3952,s3887,s3878,s3930);
  nand x1509(s3966,s5425,s5428);
  nand x1510(s4107,s4104,s132);
  or x1511(s4196,s1046,s1171,s1172,s1173);
  nor x1512(s4204,s1046,s1174,s1175);
  or x1513(s4212,s1064,s1176,s1177);
  nor x1514(s4220,s1064,s1178);
  or x1515(s4244,s1111,s1188,s1189,s1190,s1191);
  or x1516(s4252,s1128,s1192,s1193,s1194);
  or x1517(s4260,s1145,s1195,s1196);
  or x1518(s4268,s1160,s1197);
  or x1519(s4361,s1301,s1442,s1443,s1444);
  nor x1520(s4419,s1301,s1445,s1446);
  or x1521(s4467,s1382,s1472,s1473,s1474);
  or x1522(s4487,s1359,s1465,s1466,s1467,s1468);
  nor x1523(s4555,s1382,s1475,s1476);
  nor x1524(s4575,s1359,s1469,s1470,s1471);
  or x1525(s4684,s1724,s1849,s1850,s1851);
  nor x1526(s4692,s1724,s1852,s1853);
  or x1527(s4700,s1742,s1854,s1855);
  nor x1528(s4708,s1742,s1856);
  or x1529(s4732,s1789,s1866,s1867,s1868,s1869);
  or x1530(s4740,s1806,s1870,s1871,s1872);
  or x1531(s4748,s1823,s1873,s1874);
  or x1532(s4825,s1978,s2119,s2120,s2121);
  nor x1533(s4883,s1978,s2122,s2123);
  or x1534(s4928,s2059,s2149,s2150,s2151);
  or x1535(s4941,s2036,s2142,s2143,s2144,s2145);
  nor x1536(s5009,s2059,s2152,s2153);
  nor x1537(s5029,s2036,s2146,s2147,s2148);
  nand x1538(s5224,s5219,s5222);
  nand x1539(s5225,s5216,s5223);
  nand x1540(s5234,s5229,s5232);
  nand x1541(s5235,s5226,s5233);
  nand x1542(s5376,s5294,s5295);
  nand x1543(s5417,s5394,s5395);
  not x1544(s576,s1878);
  and x1545(s588,s1437,s1451);
  and x1546(s615,s1843,s1857);
  and x1547(s626,s2113,s2128);
  and x1548(s632,s1166,s1179);
  nand x1549(s1198,s4191,s4194);
  not x1550(s4195,s4191);
  not x1551(s4203,s4199);
  not x1552(s4211,s4207);
  not x1553(s4219,s4215);
  not x1554(s4227,s4223);
  nand x1555(s1217,s4231,s4234);
  not x1556(s4235,s4231);
  nand x1557(s1221,s4239,s4242);
  not x1558(s4243,s4239);
  and x1559(s1224,s1179,s4);
  not x1560(s4251,s4247);
  not x1561(s4259,s4255);
  not x1562(s4267,s4263);
  not x1563(s4275,s4271);
  not x1564(s1453,s1451);
  not x1565(s4405,s4401);
  not x1566(s4463,s4459);
  not x1567(s4541,s4537);
  not x1568(s4551,s4547);
  nand x1569(s1895,s4719,s4722);
  not x1570(s4723,s4719);
  nand x1571(s1899,s4727,s4730);
  not x1572(s4731,s4727);
  and x1573(s1902,s1857,s54);
  not x1574(s4739,s4735);
  not x1575(s4755,s4751);
  nand x1576(s1929,s4759,s4762);
  not x1577(s4763,s4759);
  not x1578(s2130,s2128);
  not x1579(s3500,s3497);
  not x1580(s3504,s3501);
  not x1581(s3508,s3505);
  not x1582(s3512,s3509);
  and x1583(s3520,s3454,s3445,s3497);
  and x1584(s3523,s3458,s3449,s3501);
  and x1585(s3526,s3477,s3468,s3505);
  and x1586(s3529,s3481,s3472,s3509);
  buf x1587(s1002,s3533);
  and x1588(s3837,s1878,s3795,s3823);
  and x1589(s3942,s3857,s3862,s3921);
  and x1590(s3945,s3853,s3866,s3925);
  and x1591(s3948,s3878,s3883,s3929);
  and x1592(s3951,s3874,s3887,s3933);
  nand x1593(s3968,s3966,s3967);
  not x1594(s4375,s4371);
  not x1595(s4385,s4381);
  not x1596(s4395,s4391);
  not x1597(s4433,s4429);
  not x1598(s4443,s4439);
  not x1599(s4453,s4449);
  not x1600(s4501,s4497);
  not x1601(s4511,s4507);
  not x1602(s4521,s4517);
  not x1603(s4531,s4527);
  not x1604(s4619,s4615);
  not x1605(s4589,s4585);
  not x1606(s4599,s4595);
  not x1607(s4609,s4605);
  not x1608(s4839,s4835);
  not x1609(s4849,s4845);
  not x1610(s4897,s4893);
  not x1611(s4907,s4903);
  not x1612(s4965,s4961);
  not x1613(s4975,s4971);
  not x1614(s4985,s4981);
  not x1615(s5073,s5069);
  not x1616(s5053,s5049);
  not x1617(s5063,s5059);
  nand x1618(s5247,s5224,s5225);
  nand x1619(s5255,s5234,s5235);
  and x1620(s590,s1437,s1458);
  and x1621(s617,s1863,s1843);
  and x1622(s620,s1185,s1166);
  and x1623(s628,s2113,s2135);
  not x1624(s3535,s3533);
  nand x1625(s1199,s4188,s4195);
  not x1626(s4202,s4196);
  nand x1627(s1204,s4196,s4203);
  not x1628(s4210,s4204);
  nand x1629(s1207,s4204,s4211);
  not x1630(s4218,s4212);
  nand x1631(s1211,s4212,s4219);
  not x1632(s4226,s4220);
  nand x1633(s1214,s4220,s4227);
  nand x1634(s1218,s4228,s4235);
  nand x1635(s1222,s4236,s4243);
  or x1636(s1225,s1185,s1224);
  not x1637(s4250,s4244);
  nand x1638(s1237,s4244,s4251);
  not x1639(s4258,s4252);
  nand x1640(s1242,s4252,s4259);
  not x1641(s4266,s4260);
  nand x1642(s1247,s4260,s4267);
  not x1643(s4274,s4268);
  nand x1644(s1252,s4268,s4275);
  not x1645(s1462,s1458);
  not x1646(s4690,s4684);
  nand x1647(s1882,s4684,s4691);
  not x1648(s4698,s4692);
  nand x1649(s1885,s4692,s4699);
  not x1650(s4706,s4700);
  nand x1651(s1889,s4700,s4707);
  not x1652(s4714,s4708);
  nand x1653(s1892,s4708,s4715);
  nand x1654(s1896,s4716,s4723);
  nand x1655(s1900,s4724,s4731);
  or x1656(s1903,s1863,s1902);
  not x1657(s4738,s4732);
  nand x1658(s1915,s4732,s4739);
  not x1659(s4746,s4740);
  nand x1660(s1920,s4740,s4747);
  not x1661(s4754,s4748);
  nand x1662(s1925,s4748,s4755);
  nand x1663(s1930,s4756,s4763);
  not x1664(s2139,s2135);
  and x1665(s3519,s3449,s3454,s3500);
  and x1666(s3522,s3445,s3458,s3504);
  and x1667(s3525,s3472,s3477,s3508);
  and x1668(s3528,s3468,s3481,s3512);
  or x1669(s3848,s3836,s3837,s3838);
  nor x1670(s3944,s3942,s3943);
  nor x1671(s3947,s3945,s3946);
  nor x1672(s3950,s3948,s3949);
  nor x1673(s3953,s3951,s3952);
  not x1674(s5421,s5417);
  buf x1675(s1004,s3968);
  and x1676(s4111,s4104,s4107);
  and x1677(s4112,s4107,s132);
  or x1678(s4351,s1448,s1481);
  not x1679(s4365,s4361);
  not x1680(s4409,s1448);
  not x1681(s4423,s4419);
  not x1682(s4471,s4467);
  nand x1683(s4472,s4467,s4470);
  or x1684(s4477,s1478,s1482);
  not x1685(s4491,s4487);
  not x1686(s4559,s4555);
  nand x1687(s4560,s4555,s4558);
  not x1688(s4565,s1478);
  not x1689(s4579,s4575);
  or x1690(s4815,s2125,s2158);
  not x1691(s4829,s4825);
  not x1692(s4873,s2125);
  not x1693(s4887,s4883);
  or x1694(s4931,s2155,s2159);
  not x1695(s4934,s4928);
  not x1696(s4945,s4941);
  not x1697(s5013,s5009);
  nand x1698(s5014,s5009,s5012);
  not x1699(s5019,s2155);
  not x1700(s5033,s5029);
  not x1701(s5382,s5376);
  nand x1702(s5385,s5376,s5383);
  or x1703(s591,s589,s590);
  or x1704(s618,s616,s617);
  or x1705(s621,s619,s620);
  or x1706(s629,s627,s628);
  not x1707(s3970,s3968);
  nand x1708(s1200,s1198,s1199);
  nand x1709(s1203,s4199,s4202);
  nand x1710(s1206,s4207,s4210);
  nand x1711(s1210,s4215,s4218);
  nand x1712(s1213,s4223,s4226);
  nand x1713(s1219,s1217,s1218);
  nand x1714(s1223,s1221,s1222);
  nand x1715(s1236,s4247,s4250);
  nand x1716(s1241,s4255,s4258);
  nand x1717(s1246,s4263,s4266);
  nand x1718(s1251,s4271,s4274);
  nand x1719(s1881,s4687,s4690);
  nand x1720(s1884,s4695,s4698);
  nand x1721(s1888,s4703,s4706);
  nand x1722(s1891,s4711,s4714);
  nand x1723(s1897,s1895,s1896);
  nand x1724(s1901,s1899,s1900);
  nand x1725(s1914,s4735,s4738);
  nand x1726(s1919,s4743,s4746);
  nand x1727(s1924,s4751,s4754);
  nand x1728(s1931,s1929,s1930);
  nor x1729(s3521,s3519,s3520);
  nor x1730(s3524,s3522,s3523);
  nor x1731(s3527,s3525,s3526);
  nor x1732(s3530,s3528,s3529);
  not x1733(s5251,s5247);
  not x1734(s5259,s5255);
  or x1735(s4113,s4111,s4112);
  nand x1736(s4473,s4464,s4471);
  nand x1737(s4561,s4552,s4559);
  nand x1738(s5015,s5006,s5013);
  nand x1739(s5384,s5379,s5382);
  nand x1740(s5406,s3947,s3944);
  nand x1741(s5414,s3953,s3950);
  and x1742(s1664,s3848,s1621,s1645);
  and x1743(s2335,s3848,s2293,s2316);
  and x1744(s718,s3848,s2430,s2454);
  not x1745(s822,s3848);
  and x1746(s855,s3848,s2488,s2512);
  nand x1747(s1205,s1203,s1204);
  nand x1748(s1208,s1206,s1207);
  nand x1749(s1212,s1210,s1211);
  nand x1750(s1215,s1213,s1214);
  not x1751(s1220,s1219);
  not x1752(s1231,s1225);
  nand x1753(s1238,s1236,s1237);
  nand x1754(s1243,s1241,s1242);
  nand x1755(s1248,s1246,s1247);
  nand x1756(s1253,s1251,s1252);
  and x1757(s1272,s1225,s1086);
  and x1758(s1483,s1462,s1453);
  nand x1759(s1883,s1881,s1882);
  nand x1760(s1886,s1884,s1885);
  nand x1761(s1890,s1888,s1889);
  nand x1762(s1893,s1891,s1892);
  not x1763(s1898,s1897);
  not x1764(s1909,s1903);
  nand x1765(s1916,s1914,s1915);
  nand x1766(s1921,s1919,s1920);
  nand x1767(s1926,s1924,s1925);
  and x1768(s1953,s1903,s1764);
  and x1769(s2160,s2139,s2130);
  not x1770(s4355,s4351);
  nand x1771(s4356,s4351,s4354);
  not x1772(s4413,s4409);
  nand x1773(s4414,s4409,s4412);
  nand x1774(s4474,s4472,s4473);
  not x1775(s4481,s4477);
  nand x1776(s4562,s4560,s4561);
  not x1777(s4569,s4565);
  not x1778(s4819,s4815);
  nand x1779(s4820,s4815,s4818);
  not x1780(s4877,s4873);
  nand x1781(s4878,s4873,s4876);
  not x1782(s4935,s4931);
  nand x1783(s4936,s4931,s4934);
  nand x1784(s5016,s5014,s5015);
  not x1785(s5023,s5019);
  nand x1786(s5244,s3524,s3521);
  nand x1787(s5252,s3530,s3527);
  nand x1788(s5409,s5384,s5385);
  not x1789(s566,s1200);
  not x1790(s577,s1931);
  and x1791(s3733,s4113,s3724,s3721);
  not x1792(s1209,s1208);
  not x1793(s1216,s1215);
  and x1794(s1257,s1225,s1205);
  and x1795(s1262,s1225,s1212);
  and x1796(s1267,s1225,s1220);
  not x1797(s1887,s1886);
  not x1798(s1894,s1893);
  and x1799(s1935,s1903,s1883);
  and x1800(s1943,s1903,s1890);
  and x1801(s1948,s1903,s1898);
  and x1802(s3779,s1200,s3737,s3765);
  and x1803(s3840,s1931,s3795,s3823);
  not x1804(s5412,s5406);
  not x1805(s5420,s5414);
  nand x1806(s3964,s5414,s5421);
  nand x1807(s4357,s4348,s4355);
  nand x1808(s4415,s4406,s4413);
  nand x1809(s4821,s4812,s4819);
  nand x1810(s4879,s4870,s4877);
  nand x1811(s4937,s4928,s4935);
  not x1812(s567,s1253);
  not x1813(s568,s1248);
  not x1814(s569,s1243);
  not x1815(s570,s1238);
  not x1816(s578,s1926);
  not x1817(s579,s1921);
  not x1818(s580,s1916);
  and x1819(s1256,s1209,s1231);
  and x1820(s1261,s1216,s1231);
  and x1821(s1266,s1223,s1231);
  and x1822(s1271,s1080,s1231);
  not x1823(s1486,s1483);
  and x1824(s1934,s1887,s1909);
  and x1825(s1942,s1894,s1909);
  and x1826(s1947,s1901,s1909);
  and x1827(s1952,s1758,s1909);
  not x1828(s2163,s2160);
  not x1829(s5250,s5244);
  nand x1830(s3537,s5244,s5251);
  not x1831(s5258,s5252);
  nand x1832(s3542,s5252,s5259);
  and x1833(s3782,s1253,s3737,s3765);
  and x1834(s3785,s1248,s3737,s3765);
  and x1835(s3788,s1243,s3737,s3765);
  or x1836(s3790,s3778,s3779,s3780);
  and x1837(s3843,s1926,s3795,s3823);
  and x1838(s3846,s1921,s3795,s3823);
  or x1839(s3849,s3839,s3840,s3841);
  nand x1840(s3960,s5409,s5412);
  not x1841(s5413,s5409);
  nand x1842(s3963,s5417,s5420);
  and x1843(s4010,s1238,s3972,s3998);
  and x1844(s4068,s1916,s4030,s4056);
  nand x1845(s4358,s4356,s4357);
  nand x1846(s4416,s4414,s4415);
  not x1847(s4480,s4474);
  nand x1848(s4483,s4474,s4481);
  not x1849(s4568,s4562);
  nand x1850(s4571,s4562,s4569);
  nand x1851(s4822,s4820,s4821);
  nand x1852(s4880,s4878,s4879);
  nand x1853(s4938,s4936,s4937);
  not x1854(s5022,s5016);
  nand x1855(s5025,s5016,s5023);
  or x1856(s1258,s1256,s1257);
  or x1857(s1263,s1261,s1262);
  or x1858(s1268,s1266,s1267);
  or x1859(s1273,s1271,s1272);
  or x1860(s1936,s1934,s1935);
  or x1861(s1944,s1942,s1943);
  or x1862(s1949,s1947,s1948);
  or x1863(s1954,s1952,s1953);
  nand x1864(s3536,s5247,s5250);
  nand x1865(s3541,s5255,s5258);
  or x1866(s3791,s3781,s3782,s3783);
  or x1867(s3792,s3784,s3785,s3786);
  or x1868(s3793,s3787,s3788,s3789);
  or x1869(s3850,s3842,s3843,s3844);
  or x1870(s3851,s3845,s3846,s3847);
  nand x1871(s3961,s5406,s5413);
  nand x1872(s3965,s3963,s3964);
  or x1873(s4024,s4009,s4010,s4011);
  or x1874(s4082,s4067,s4068,s4069);
  nand x1875(s4482,s4477,s4480);
  nand x1876(s4570,s4565,s4568);
  nand x1877(s5024,s5019,s5022);
  and x1878(s1666,s3790,s1609,s1645);
  and x1879(s1670,s3849,s1621,s1645);
  and x1880(s2337,s3790,s2281,s2316);
  and x1881(s2341,s3849,s2293,s2316);
  and x1882(s719,s3790,s2418,s2454);
  and x1883(s758,s3849,s2430,s2454);
  and x1884(s798,s3849,s2488,s2512);
  not x1885(s838,s3849);
  and x1886(s856,s3790,s2476,s2512);
  not x1887(s861,s3790);
  nand x1888(s3538,s3536,s3537);
  nand x1889(s3543,s3541,s3542);
  nand x1890(s3962,s3960,s3961);
  not x1891(s4364,s4358);
  nand x1892(s4367,s4358,s4365);
  not x1893(s4422,s4416);
  nand x1894(s4425,s4416,s4423);
  nand x1895(s4484,s4482,s4483);
  nand x1896(s4572,s4570,s4571);
  not x1897(s4828,s4822);
  nand x1898(s4831,s4822,s4829);
  not x1899(s4886,s4880);
  nand x1900(s4889,s4880,s4887);
  not x1901(s4944,s4938);
  nand x1902(s4947,s4938,s4945);
  nand x1903(s5026,s5024,s5025);
  not x1904(s571,s1273);
  not x1905(s572,s1268);
  not x1906(s573,s1263);
  not x1907(s574,s1258);
  not x1908(s581,s1954);
  not x1909(s582,s1949);
  not x1910(s583,s1944);
  not x1911(s584,s1936);
  not x1912(s623,s1936);
  and x1913(s1576,s4082,s1540,s1564);
  and x1914(s1578,s4024,s1528,s1564);
  or x1915(s659,s1664,s1666,s1667,s1668);
  and x1916(s1672,s3791,s1609,s1645);
  and x1917(s1676,s3850,s1621,s1645);
  and x1918(s1678,s3792,s1609,s1645);
  and x1919(s1682,s3851,s1621,s1645);
  and x1920(s1684,s3793,s1609,s1645);
  and x1921(s2250,s4082,s2215,s2238);
  and x1922(s2252,s4024,s2203,s2238);
  or x1923(s691,s2335,s2337,s2338,s2339);
  and x1924(s2343,s3791,s2281,s2316);
  and x1925(s2347,s3850,s2293,s2316);
  and x1926(s2349,s3792,s2281,s2316);
  and x1927(s2353,s3851,s2293,s2316);
  and x1928(s2355,s3793,s2281,s2316);
  or x1929(s722,s718,s719,s720,s721);
  and x1930(s743,s4082,s3570,s3594);
  and x1931(s744,s4024,s3558,s3594);
  and x1932(s748,s3851,s2430,s2454);
  and x1933(s749,s3793,s2418,s2454);
  and x1934(s753,s3850,s2430,s2454);
  and x1935(s754,s3792,s2418,s2454);
  and x1936(s759,s3791,s2418,s2454);
  and x1937(s783,s4082,s3672,s3696);
  and x1938(s784,s4024,s3660,s3696);
  and x1939(s788,s3851,s2488,s2512);
  and x1940(s789,s3793,s2476,s2512);
  and x1941(s793,s3850,s2488,s2512);
  and x1942(s794,s3792,s2476,s2512);
  and x1943(s799,s3791,s2476,s2512);
  and x1944(s3735,s1936,s3724,s3717);
  not x1945(s832,s4082);
  not x1946(s834,s3851);
  not x1947(s836,s3850);
  not x1948(s3835,s3965);
  or x1949(s859,s855,s856,s857,s858);
  not x1950(s871,s4024);
  not x1951(s873,s3793);
  not x1952(s875,s3792);
  not x1953(s877,s3791);
  buf x1954(s998,s3538);
  buf x1955(s1000,s3543);
  and x1956(s3651,s3965,s3632);
  and x1957(s4013,s1273,s3972,s3998);
  and x1958(s4016,s1268,s3972,s3998);
  and x1959(s4019,s1263,s3972,s3998);
  and x1960(s4022,s1258,s3972,s3998);
  and x1961(s4071,s1954,s4030,s4056);
  and x1962(s4074,s1949,s4030,s4056);
  and x1963(s4077,s1944,s4030,s4056);
  and x1964(s4080,s1936,s4030,s4056);
  nand x1965(s4096,s4113,s1936);
  nand x1966(s4366,s4361,s4364);
  nand x1967(s4424,s4419,s4422);
  nand x1968(s4830,s4825,s4828);
  nand x1969(s4888,s4883,s4886);
  nand x1970(s4946,s4941,s4944);
  and x1971(s575,s566,s567,s568,s569,s570,s571,s572,s573,s574);
  and x1972(s585,s576,s577,s578,s579,s580,s581,s582,s583,s584);
  or x1973(s640,s1576,s1578,s1579,s1580);
  and x1974(s661,s659,s1606);
  or x1975(s662,s1670,s1672,s1673,s1674);
  or x1976(s665,s1676,s1678,s1679,s1680);
  or x1977(s668,s1682,s1684,s1685,s1686);
  or x1978(s674,s2250,s2252,s2253,s2254);
  and x1979(s693,s691,s2279);
  or x1980(s694,s2341,s2343,s2344,s2345);
  or x1981(s697,s2347,s2349,s2350,s2351);
  or x1982(s700,s2353,s2355,s2356,s2357);
  or x1983(s747,s743,s744,s745,s746);
  or x1984(s752,s748,s749,s750,s751);
  or x1985(s757,s753,s754,s755,s756);
  or x1986(s762,s758,s759,s760,s761);
  or x1987(s787,s783,s784,s785,s786);
  or x1988(s792,s788,s789,s790,s791);
  or x1989(s797,s793,s794,s795,s796);
  or x1990(s802,s798,s799,s800,s801);
  or x1991(s817,s3731,s3733,s3734,s3735);
  and x1992(s839,s3835,s3803,s3823);
  not x1993(s3540,s3538);
  not x1994(s3545,s3543);
  not x1995(s3777,s3962);
  and x1996(s3648,s3962,s3632);
  or x1997(s4025,s4012,s4013,s4014);
  or x1998(s4026,s4015,s4016,s4017);
  or x1999(s4027,s4018,s4019,s4020);
  or x2000(s4028,s4021,s4022,s4023);
  or x2001(s4083,s4070,s4071,s4072);
  or x2002(s4084,s4073,s4074,s4075);
  or x2003(s4085,s4076,s4077,s4078);
  or x2004(s4086,s4079,s4080,s4081);
  nand x2005(s4368,s4366,s4367);
  nand x2006(s4426,s4424,s4425);
  not x2007(s4490,s4484);
  nand x2008(s4493,s4484,s4491);
  not x2009(s4578,s4572);
  nand x2010(s4581,s4572,s4579);
  nand x2011(s4832,s4830,s4831);
  nand x2012(s4890,s4888,s4889);
  nand x2013(s4948,s4946,s4947);
  not x2014(s5032,s5026);
  nand x2015(s5035,s5026,s5033);
  and x2016(s642,s640,s1526);
  and x2017(s664,s662,s1606);
  and x2018(s667,s665,s1606);
  and x2019(s670,s668,s1606);
  and x2020(s676,s674,s2202);
  and x2021(s696,s694,s2279);
  and x2022(s699,s697,s2279);
  and x2023(s702,s700,s2279);
  and x2024(s811,s4113,s4096);
  and x2025(s812,s4096,s1936);
  and x2026(s818,s816,s817);
  and x2027(s853,s562,s3540,s3545,s3535,s3970);
  and x2028(s878,s3777,s3745,s3765);
  nand x2029(s4492,s4487,s4490);
  nand x2030(s4580,s4575,s4578);
  nand x2031(s5034,s5029,s5032);
  and x2032(s1582,s4083,s1540,s1564);
  and x2033(s1584,s4025,s1528,s1564);
  and x2034(s1588,s4084,s1540,s1564);
  and x2035(s1590,s4026,s1528,s1564);
  and x2036(s1594,s4085,s1540,s1564);
  and x2037(s1596,s4027,s1528,s1564);
  and x2038(s1600,s4086,s1540,s1564);
  and x2039(s1602,s4028,s1528,s1564);
  and x2040(s2256,s4083,s2215,s2238);
  and x2041(s2258,s4025,s2203,s2238);
  and x2042(s2262,s4084,s2215,s2238);
  and x2043(s2264,s4026,s2203,s2238);
  and x2044(s2268,s4085,s2215,s2238);
  and x2045(s2270,s4027,s2203,s2238);
  and x2046(s2274,s4086,s2215,s2238);
  and x2047(s2276,s4028,s2203,s2238);
  and x2048(s708,s4086,s3672,s3696);
  and x2049(s709,s4028,s3660,s3696);
  and x2050(s723,s4086,s3570,s3594);
  and x2051(s724,s4028,s3558,s3594);
  and x2052(s728,s4085,s3570,s3594);
  and x2053(s729,s4027,s3558,s3594);
  and x2054(s733,s4084,s3570,s3594);
  and x2055(s734,s4026,s3558,s3594);
  and x2056(s738,s4083,s3570,s3594);
  and x2057(s739,s4025,s3558,s3594);
  and x2058(s768,s4085,s3672,s3696);
  and x2059(s769,s4027,s3660,s3696);
  and x2060(s773,s4084,s3672,s3696);
  and x2061(s774,s4026,s3660,s3696);
  and x2062(s778,s4083,s3672,s3696);
  and x2063(s779,s4025,s3660,s3696);
  or x2064(s813,s811,s812);
  not x2065(s824,s4086);
  not x2066(s826,s4085);
  not x2067(s828,s4084);
  not x2068(s830,s4083);
  and x2069(s854,s852,s853,s245);
  not x2070(s863,s4028);
  not x2071(s865,s4027);
  not x2072(s867,s4026);
  not x2073(s869,s4025);
  not x2074(s4374,s4368);
  nand x2075(s4377,s4368,s4375);
  not x2076(s4432,s4426);
  nand x2077(s4435,s4426,s4433);
  nand x2078(s4494,s4492,s4493);
  nand x2079(s4582,s4580,s4581);
  not x2080(s4838,s4832);
  nand x2081(s4841,s4832,s4839);
  not x2082(s4896,s4890);
  nand x2083(s4899,s4890,s4897);
  not x2084(s4954,s4948);
  nand x2085(s4957,s4948,s4955);
  nand x2086(s5036,s5034,s5035);
  or x2087(s643,s1582,s1584,s1585,s1586);
  or x2088(s646,s1588,s1590,s1591,s1592);
  or x2089(s649,s1594,s1596,s1597,s1598);
  or x2090(s652,s1600,s1602,s1603,s1604);
  or x2091(s677,s2256,s2258,s2259,s2260);
  or x2092(s680,s2262,s2264,s2265,s2266);
  or x2093(s683,s2268,s2270,s2271,s2272);
  or x2094(s686,s2274,s2276,s2277,s2278);
  or x2095(s712,s708,s709,s710,s711);
  or x2096(s727,s723,s724,s725,s726);
  or x2097(s732,s728,s729,s730,s731);
  or x2098(s737,s733,s734,s735,s736);
  or x2099(s742,s738,s739,s740,s741);
  or x2100(s772,s768,s769,s770,s771);
  or x2101(s777,s773,s774,s775,s776);
  or x2102(s782,s778,s779,s780,s781);
  nand x2103(s4376,s4371,s4374);
  nand x2104(s4434,s4429,s4432);
  nand x2105(s4840,s4835,s4838);
  nand x2106(s4898,s4893,s4896);
  nand x2107(s4956,s4951,s4954);
  and x2108(s645,s643,s1526);
  and x2109(s648,s646,s1526);
  and x2110(s651,s649,s1526);
  and x2111(s654,s652,s1526);
  and x2112(s679,s677,s2202);
  and x2113(s682,s680,s2202);
  and x2114(s685,s683,s2202);
  and x2115(s688,s686,s2202);
  nand x2116(s4378,s4376,s4377);
  nand x2117(s4436,s4434,s4435);
  not x2118(s4500,s4494);
  nand x2119(s4503,s4494,s4501);
  not x2120(s4588,s4582);
  nand x2121(s4591,s4582,s4589);
  nand x2122(s4842,s4840,s4841);
  nand x2123(s4900,s4898,s4899);
  nand x2124(s4958,s4956,s4957);
  not x2125(s5042,s5036);
  nand x2126(s5045,s5036,s5043);
  nand x2127(s4502,s4497,s4500);
  nand x2128(s4590,s4585,s4588);
  nand x2129(s5044,s5039,s5042);
  not x2130(s4384,s4378);
  nand x2131(s4387,s4378,s4385);
  not x2132(s4442,s4436);
  nand x2133(s4445,s4436,s4443);
  nand x2134(s4504,s4502,s4503);
  nand x2135(s4592,s4590,s4591);
  not x2136(s4848,s4842);
  nand x2137(s4851,s4842,s4849);
  not x2138(s4906,s4900);
  nand x2139(s4909,s4900,s4907);
  not x2140(s4964,s4958);
  nand x2141(s4967,s4958,s4965);
  nand x2142(s5046,s5044,s5045);
  nand x2143(s4386,s4381,s4384);
  nand x2144(s4444,s4439,s4442);
  nand x2145(s4850,s4845,s4848);
  nand x2146(s4908,s4903,s4906);
  nand x2147(s4966,s4961,s4964);
  nand x2148(s4388,s4386,s4387);
  nand x2149(s4446,s4444,s4445);
  not x2150(s4510,s4504);
  nand x2151(s4513,s4504,s4511);
  not x2152(s4598,s4592);
  nand x2153(s4601,s4592,s4599);
  nand x2154(s4852,s4850,s4851);
  nand x2155(s4910,s4908,s4909);
  nand x2156(s4968,s4966,s4967);
  not x2157(s5052,s5046);
  nand x2158(s5055,s5046,s5053);
  nand x2159(s4512,s4507,s4510);
  nand x2160(s4600,s4595,s4598);
  nand x2161(s5054,s5049,s5052);
  not x2162(s4394,s4388);
  nand x2163(s4397,s4388,s4395);
  not x2164(s4452,s4446);
  nand x2165(s4455,s4446,s4453);
  nand x2166(s4514,s4512,s4513);
  nand x2167(s4602,s4600,s4601);
  not x2168(s4858,s4852);
  nand x2169(s4861,s4852,s4859);
  not x2170(s4916,s4910);
  nand x2171(s4919,s4910,s4917);
  not x2172(s4974,s4968);
  nand x2173(s4977,s4968,s4975);
  nand x2174(s5056,s5054,s5055);
  nand x2175(s4396,s4391,s4394);
  nand x2176(s4454,s4449,s4452);
  nand x2177(s4860,s4855,s4858);
  nand x2178(s4918,s4913,s4916);
  nand x2179(s4976,s4971,s4974);
  nand x2180(s4398,s4396,s4397);
  nand x2181(s4456,s4454,s4455);
  not x2182(s4520,s4514);
  nand x2183(s4523,s4514,s4521);
  not x2184(s4608,s4602);
  nand x2185(s4611,s4602,s4609);
  nand x2186(s4862,s4860,s4861);
  nand x2187(s4920,s4918,s4919);
  nand x2188(s4978,s4976,s4977);
  not x2189(s5062,s5056);
  nand x2190(s5065,s5056,s5063);
  nand x2191(s4522,s4517,s4520);
  nand x2192(s4610,s4605,s4608);
  nand x2193(s5064,s5059,s5062);
  not x2194(s4404,s4398);
  nand x2195(s1488,s4398,s4405);
  not x2196(s4462,s4456);
  nand x2197(s1493,s4456,s4463);
  not x2198(s4868,s4862);
  nand x2199(s2165,s4862,s4869);
  not x2200(s4926,s4920);
  nand x2201(s2170,s4920,s4927);
  nand x2202(s4524,s4522,s4523);
  nand x2203(s4612,s4610,s4611);
  not x2204(s4984,s4978);
  nand x2205(s4987,s4978,s4985);
  nand x2206(s5066,s5064,s5065);
  nand x2207(s1487,s4401,s4404);
  nand x2208(s1492,s4459,s4462);
  nand x2209(s2164,s4865,s4868);
  nand x2210(s2169,s4923,s4926);
  nand x2211(s4986,s4981,s4984);
  nand x2212(s1489,s1487,s1488);
  nand x2213(s1494,s1492,s1493);
  nand x2214(s2166,s2164,s2165);
  nand x2215(s2171,s2169,s2170);
  not x2216(s4530,s4524);
  nand x2217(s4533,s4524,s4531);
  not x2218(s4618,s4612);
  nand x2219(s4543,s4612,s4619);
  nand x2220(s4988,s4986,s4987);
  not x2221(s5072,s5066);
  nand x2222(s4997,s5066,s5073);
  nand x2223(s4532,s4527,s4530);
  nand x2224(s4542,s4615,s4618);
  nand x2225(s4996,s5069,s5072);
  and x2226(s1513,s1494,s1462,s1502);
  and x2227(s1514,s1489,s1458,s1502);
  and x2228(s1515,s1494,s1483,s1497);
  and x2229(s1516,s1489,s1486,s1497);
  not x2230(s4994,s4988);
  nand x2231(s2184,s4988,s4995);
  and x2232(s2190,s2171,s2139,s2179);
  and x2233(s2191,s2166,s2135,s2179);
  and x2234(s2192,s2171,s2160,s2174);
  and x2235(s2193,s2166,s2163,s2174);
  nand x2236(s4534,s4532,s4533);
  nand x2237(s4544,s4542,s4543);
  nand x2238(s4998,s4996,s4997);
  nand x2239(s2183,s4991,s4994);
  or x2240(s4620,s1513,s1514,s1515,s1516);
  or x2241(s5074,s2190,s2191,s2192,s2193);
  not x2242(s4540,s4534);
  nand x2243(s1507,s4534,s4541);
  not x2244(s4550,s4544);
  nand x2245(s1510,s4544,s4551);
  nand x2246(s2185,s2183,s2184);
  not x2247(s5004,s4998);
  nand x2248(s2187,s4998,s5005);
  nand x2249(s1506,s4537,s4540);
  nand x2250(s1509,s4547,s4550);
  not x2251(s4626,s4620);
  nand x2252(s2186,s5001,s5004);
  and x2253(s2195,s2174,s2185);
  not x2254(s5080,s5074);
  nand x2255(s1508,s1506,s1507);
  nand x2256(s1511,s1509,s1510);
  nand x2257(s2188,s2186,s2187);
  not x2258(s1512,s1511);
  and x2259(s1518,s1497,s1508);
  not x2260(s2189,s2188);
  and x2261(s1517,s1512,s1502);
  and x2262(s2194,s2189,s2179);
  or x2263(s4623,s1517,s1518);
  or x2264(s5077,s2194,s2195);
  nand x2265(s1519,s4623,s4626);
  not x2266(s4627,s4623);
  nand x2267(s2196,s5077,s5080);
  not x2268(s5081,s5077);
  nand x2269(s1520,s4620,s4627);
  nand x2270(s2197,s5074,s5081);
  nand x2271(s1521,s1519,s1520);
  nand x2272(s2198,s2196,s2197);
  and x2273(s840,s2198,s3795,s3823);
  and x2274(s879,s1521,s3737,s3765);
  not x2275(s1524,s1521);
  not x2276(s2201,s2198);
  or x2277(s843,s839,s840,s841,s842);
  or x2278(s882,s878,s879,s880,s881);
  and x2279(s3649,s1524,s3628);
  and x2280(s3652,s2201,s3628);
  or x2281(s3657,s3648,s3649);
  or x2282(s3658,s3651,s3652);
  and x2283(s3636,s3657,s3622);
  and x2284(s3639,s3658,s3622);
  and x2285(s3642,s3657,s3622);
  and x2286(s3645,s3658,s3622);
  or x2287(s3653,s3636,s3637);
  or x2288(s3654,s3639,s3640);
  or x2289(s3655,s3642,s3643);
  or x2290(s3656,s3645,s3646);
  and x2291(s763,s3656,s2430,s2454);
  and x2292(s764,s3655,s2418,s2454);
  and x2293(s803,s3656,s2488,s2512);
  and x2294(s804,s3655,s2476,s2512);
  and x2295(s1657,s3654,s1621,s1645);
  and x2296(s1659,s3653,s1609,s1645);
  and x2297(s2328,s3654,s2293,s2316);
  and x2298(s2330,s3653,s2281,s2316);
  or x2299(s1662,s1657,s1659,s1660,s1661);
  or x2300(s2333,s2328,s2330,s2331,s2332);
  or x2301(s767,s763,s764,s765,s766);
  or x2302(s807,s803,s804,s805,s806);
  and x2303(s657,s1662,s1606);
  and x2304(s689,s2333,s2279);
  not x2305(s658,s657);
  not x2306(s690,s689);

endmodule
