module c6288(s545gat,s1581gat,s1901gat,s2223gat,s2548gat,s2877gat,s3211gat,s3552gat,s3895gat,s4241gat,s4591gat,s4946gat,s5308gat,s5672gat,s5971gat,s6123gat,s6150gat,s6160gat,s6170gat,s6180gat,s6190gat,s6200gat,s6210gat,s6220gat,s6230gat,s6240gat,s6250gat,s6260gat,s6270gat,s6280gat,s6287gat,s6288gat,s1gat,s18gat,s35gat,s52gat,s69gat,s86gat,s103gat,s120gat,s137gat,s154gat,s171gat,s188gat,s205gat,s222gat,s239gat,s256gat,s273gat,s290gat,s307gat,s324gat,s341gat,s358gat,s375gat,s392gat,s409gat,s426gat,s443gat,s460gat,s477gat,s494gat,s511gat,s528gat);

  output s545gat;
  output s1581gat;
  output s1901gat;
  output s2223gat;
  output s2548gat;
  output s2877gat;
  output s3211gat;
  output s3552gat;
  output s3895gat;
  output s4241gat;
  output s4591gat;
  output s4946gat;
  output s5308gat;
  output s5672gat;
  output s5971gat;
  output s6123gat;
  output s6150gat;
  output s6160gat;
  output s6170gat;
  output s6180gat;
  output s6190gat;
  output s6200gat;
  output s6210gat;
  output s6220gat;
  output s6230gat;
  output s6240gat;
  output s6250gat;
  output s6260gat;
  output s6270gat;
  output s6280gat;
  output s6287gat;
  output s6288gat;
  input s1gat;
  input s18gat;
  input s35gat;
  input s52gat;
  input s69gat;
  input s86gat;
  input s103gat;
  input s120gat;
  input s137gat;
  input s154gat;
  input s171gat;
  input s188gat;
  input s205gat;
  input s222gat;
  input s239gat;
  input s256gat;
  input s273gat;
  input s290gat;
  input s307gat;
  input s324gat;
  input s341gat;
  input s358gat;
  input s375gat;
  input s392gat;
  input s409gat;
  input s426gat;
  input s443gat;
  input s460gat;
  input s477gat;
  input s494gat;
  input s511gat;
  input s528gat;

  and x0(s545gat,s1gat,s273gat);
  and x1(s546gat,s1gat,s290gat);
  and x2(s549gat,s1gat,s307gat);
  and x3(s552gat,s1gat,s324gat);
  and x4(s555gat,s1gat,s341gat);
  and x5(s558gat,s1gat,s358gat);
  and x6(s561gat,s1gat,s375gat);
  and x7(s564gat,s1gat,s392gat);
  and x8(s567gat,s1gat,s409gat);
  and x9(s570gat,s1gat,s426gat);
  and x10(s573gat,s1gat,s443gat);
  and x11(s576gat,s1gat,s460gat);
  and x12(s579gat,s1gat,s477gat);
  and x13(s582gat,s1gat,s494gat);
  and x14(s585gat,s1gat,s511gat);
  and x15(s588gat,s1gat,s528gat);
  and x16(s591gat,s18gat,s273gat);
  and x17(s594gat,s18gat,s290gat);
  and x18(s597gat,s18gat,s307gat);
  and x19(s600gat,s18gat,s324gat);
  and x20(s603gat,s18gat,s341gat);
  and x21(s606gat,s18gat,s358gat);
  and x22(s609gat,s18gat,s375gat);
  and x23(s612gat,s18gat,s392gat);
  and x24(s615gat,s18gat,s409gat);
  and x25(s618gat,s18gat,s426gat);
  and x26(s621gat,s18gat,s443gat);
  and x27(s624gat,s18gat,s460gat);
  and x28(s627gat,s18gat,s477gat);
  and x29(s630gat,s18gat,s494gat);
  and x30(s633gat,s18gat,s511gat);
  and x31(s636gat,s18gat,s528gat);
  and x32(s639gat,s35gat,s273gat);
  and x33(s642gat,s35gat,s290gat);
  and x34(s645gat,s35gat,s307gat);
  and x35(s648gat,s35gat,s324gat);
  and x36(s651gat,s35gat,s341gat);
  and x37(s654gat,s35gat,s358gat);
  and x38(s657gat,s35gat,s375gat);
  and x39(s660gat,s35gat,s392gat);
  and x40(s663gat,s35gat,s409gat);
  and x41(s666gat,s35gat,s426gat);
  and x42(s669gat,s35gat,s443gat);
  and x43(s672gat,s35gat,s460gat);
  and x44(s675gat,s35gat,s477gat);
  and x45(s678gat,s35gat,s494gat);
  and x46(s681gat,s35gat,s511gat);
  and x47(s684gat,s35gat,s528gat);
  and x48(s687gat,s52gat,s273gat);
  and x49(s690gat,s52gat,s290gat);
  and x50(s693gat,s52gat,s307gat);
  and x51(s696gat,s52gat,s324gat);
  and x52(s699gat,s52gat,s341gat);
  and x53(s702gat,s52gat,s358gat);
  and x54(s705gat,s52gat,s375gat);
  and x55(s708gat,s52gat,s392gat);
  and x56(s711gat,s52gat,s409gat);
  and x57(s714gat,s52gat,s426gat);
  and x58(s717gat,s52gat,s443gat);
  and x59(s720gat,s52gat,s460gat);
  and x60(s723gat,s52gat,s477gat);
  and x61(s726gat,s52gat,s494gat);
  and x62(s729gat,s52gat,s511gat);
  and x63(s732gat,s52gat,s528gat);
  and x64(s735gat,s69gat,s273gat);
  and x65(s738gat,s69gat,s290gat);
  and x66(s741gat,s69gat,s307gat);
  and x67(s744gat,s69gat,s324gat);
  and x68(s747gat,s69gat,s341gat);
  and x69(s750gat,s69gat,s358gat);
  and x70(s753gat,s69gat,s375gat);
  and x71(s756gat,s69gat,s392gat);
  and x72(s759gat,s69gat,s409gat);
  and x73(s762gat,s69gat,s426gat);
  and x74(s765gat,s69gat,s443gat);
  and x75(s768gat,s69gat,s460gat);
  and x76(s771gat,s69gat,s477gat);
  and x77(s774gat,s69gat,s494gat);
  and x78(s777gat,s69gat,s511gat);
  and x79(s780gat,s69gat,s528gat);
  and x80(s783gat,s86gat,s273gat);
  and x81(s786gat,s86gat,s290gat);
  and x82(s789gat,s86gat,s307gat);
  and x83(s792gat,s86gat,s324gat);
  and x84(s795gat,s86gat,s341gat);
  and x85(s798gat,s86gat,s358gat);
  and x86(s801gat,s86gat,s375gat);
  and x87(s804gat,s86gat,s392gat);
  and x88(s807gat,s86gat,s409gat);
  and x89(s810gat,s86gat,s426gat);
  and x90(s813gat,s86gat,s443gat);
  and x91(s816gat,s86gat,s460gat);
  and x92(s819gat,s86gat,s477gat);
  and x93(s822gat,s86gat,s494gat);
  and x94(s825gat,s86gat,s511gat);
  and x95(s828gat,s86gat,s528gat);
  and x96(s831gat,s103gat,s273gat);
  and x97(s834gat,s103gat,s290gat);
  and x98(s837gat,s103gat,s307gat);
  and x99(s840gat,s103gat,s324gat);
  and x100(s843gat,s103gat,s341gat);
  and x101(s846gat,s103gat,s358gat);
  and x102(s849gat,s103gat,s375gat);
  and x103(s852gat,s103gat,s392gat);
  and x104(s855gat,s103gat,s409gat);
  and x105(s858gat,s103gat,s426gat);
  and x106(s861gat,s103gat,s443gat);
  and x107(s864gat,s103gat,s460gat);
  and x108(s867gat,s103gat,s477gat);
  and x109(s870gat,s103gat,s494gat);
  and x110(s873gat,s103gat,s511gat);
  and x111(s876gat,s103gat,s528gat);
  and x112(s879gat,s120gat,s273gat);
  and x113(s882gat,s120gat,s290gat);
  and x114(s885gat,s120gat,s307gat);
  and x115(s888gat,s120gat,s324gat);
  and x116(s891gat,s120gat,s341gat);
  and x117(s894gat,s120gat,s358gat);
  and x118(s897gat,s120gat,s375gat);
  and x119(s900gat,s120gat,s392gat);
  and x120(s903gat,s120gat,s409gat);
  and x121(s906gat,s120gat,s426gat);
  and x122(s909gat,s120gat,s443gat);
  and x123(s912gat,s120gat,s460gat);
  and x124(s915gat,s120gat,s477gat);
  and x125(s918gat,s120gat,s494gat);
  and x126(s921gat,s120gat,s511gat);
  and x127(s924gat,s120gat,s528gat);
  and x128(s927gat,s137gat,s273gat);
  and x129(s930gat,s137gat,s290gat);
  and x130(s933gat,s137gat,s307gat);
  and x131(s936gat,s137gat,s324gat);
  and x132(s939gat,s137gat,s341gat);
  and x133(s942gat,s137gat,s358gat);
  and x134(s945gat,s137gat,s375gat);
  and x135(s948gat,s137gat,s392gat);
  and x136(s951gat,s137gat,s409gat);
  and x137(s954gat,s137gat,s426gat);
  and x138(s957gat,s137gat,s443gat);
  and x139(s960gat,s137gat,s460gat);
  and x140(s963gat,s137gat,s477gat);
  and x141(s966gat,s137gat,s494gat);
  and x142(s969gat,s137gat,s511gat);
  and x143(s972gat,s137gat,s528gat);
  and x144(s975gat,s154gat,s273gat);
  and x145(s978gat,s154gat,s290gat);
  and x146(s981gat,s154gat,s307gat);
  and x147(s984gat,s154gat,s324gat);
  and x148(s987gat,s154gat,s341gat);
  and x149(s990gat,s154gat,s358gat);
  and x150(s993gat,s154gat,s375gat);
  and x151(s996gat,s154gat,s392gat);
  and x152(s999gat,s154gat,s409gat);
  and x153(s1002gat,s154gat,s426gat);
  and x154(s1005gat,s154gat,s443gat);
  and x155(s1008gat,s154gat,s460gat);
  and x156(s1011gat,s154gat,s477gat);
  and x157(s1014gat,s154gat,s494gat);
  and x158(s1017gat,s154gat,s511gat);
  and x159(s1020gat,s154gat,s528gat);
  and x160(s1023gat,s171gat,s273gat);
  and x161(s1026gat,s171gat,s290gat);
  and x162(s1029gat,s171gat,s307gat);
  and x163(s1032gat,s171gat,s324gat);
  and x164(s1035gat,s171gat,s341gat);
  and x165(s1038gat,s171gat,s358gat);
  and x166(s1041gat,s171gat,s375gat);
  and x167(s1044gat,s171gat,s392gat);
  and x168(s1047gat,s171gat,s409gat);
  and x169(s1050gat,s171gat,s426gat);
  and x170(s1053gat,s171gat,s443gat);
  and x171(s1056gat,s171gat,s460gat);
  and x172(s1059gat,s171gat,s477gat);
  and x173(s1062gat,s171gat,s494gat);
  and x174(s1065gat,s171gat,s511gat);
  and x175(s1068gat,s171gat,s528gat);
  and x176(s1071gat,s188gat,s273gat);
  and x177(s1074gat,s188gat,s290gat);
  and x178(s1077gat,s188gat,s307gat);
  and x179(s1080gat,s188gat,s324gat);
  and x180(s1083gat,s188gat,s341gat);
  and x181(s1086gat,s188gat,s358gat);
  and x182(s1089gat,s188gat,s375gat);
  and x183(s1092gat,s188gat,s392gat);
  and x184(s1095gat,s188gat,s409gat);
  and x185(s1098gat,s188gat,s426gat);
  and x186(s1101gat,s188gat,s443gat);
  and x187(s1104gat,s188gat,s460gat);
  and x188(s1107gat,s188gat,s477gat);
  and x189(s1110gat,s188gat,s494gat);
  and x190(s1113gat,s188gat,s511gat);
  and x191(s1116gat,s188gat,s528gat);
  and x192(s1119gat,s205gat,s273gat);
  and x193(s1122gat,s205gat,s290gat);
  and x194(s1125gat,s205gat,s307gat);
  and x195(s1128gat,s205gat,s324gat);
  and x196(s1131gat,s205gat,s341gat);
  and x197(s1134gat,s205gat,s358gat);
  and x198(s1137gat,s205gat,s375gat);
  and x199(s1140gat,s205gat,s392gat);
  and x200(s1143gat,s205gat,s409gat);
  and x201(s1146gat,s205gat,s426gat);
  and x202(s1149gat,s205gat,s443gat);
  and x203(s1152gat,s205gat,s460gat);
  and x204(s1155gat,s205gat,s477gat);
  and x205(s1158gat,s205gat,s494gat);
  and x206(s1161gat,s205gat,s511gat);
  and x207(s1164gat,s205gat,s528gat);
  and x208(s1167gat,s222gat,s273gat);
  and x209(s1170gat,s222gat,s290gat);
  and x210(s1173gat,s222gat,s307gat);
  and x211(s1176gat,s222gat,s324gat);
  and x212(s1179gat,s222gat,s341gat);
  and x213(s1182gat,s222gat,s358gat);
  and x214(s1185gat,s222gat,s375gat);
  and x215(s1188gat,s222gat,s392gat);
  and x216(s1191gat,s222gat,s409gat);
  and x217(s1194gat,s222gat,s426gat);
  and x218(s1197gat,s222gat,s443gat);
  and x219(s1200gat,s222gat,s460gat);
  and x220(s1203gat,s222gat,s477gat);
  and x221(s1206gat,s222gat,s494gat);
  and x222(s1209gat,s222gat,s511gat);
  and x223(s1212gat,s222gat,s528gat);
  and x224(s1215gat,s239gat,s273gat);
  and x225(s1218gat,s239gat,s290gat);
  and x226(s1221gat,s239gat,s307gat);
  and x227(s1224gat,s239gat,s324gat);
  and x228(s1227gat,s239gat,s341gat);
  and x229(s1230gat,s239gat,s358gat);
  and x230(s1233gat,s239gat,s375gat);
  and x231(s1236gat,s239gat,s392gat);
  and x232(s1239gat,s239gat,s409gat);
  and x233(s1242gat,s239gat,s426gat);
  and x234(s1245gat,s239gat,s443gat);
  and x235(s1248gat,s239gat,s460gat);
  and x236(s1251gat,s239gat,s477gat);
  and x237(s1254gat,s239gat,s494gat);
  and x238(s1257gat,s239gat,s511gat);
  and x239(s1260gat,s239gat,s528gat);
  and x240(s1263gat,s256gat,s273gat);
  and x241(s1266gat,s256gat,s290gat);
  and x242(s1269gat,s256gat,s307gat);
  and x243(s1272gat,s256gat,s324gat);
  and x244(s1275gat,s256gat,s341gat);
  and x245(s1278gat,s256gat,s358gat);
  and x246(s1281gat,s256gat,s375gat);
  and x247(s1284gat,s256gat,s392gat);
  and x248(s1287gat,s256gat,s409gat);
  and x249(s1290gat,s256gat,s426gat);
  and x250(s1293gat,s256gat,s443gat);
  and x251(s1296gat,s256gat,s460gat);
  and x252(s1299gat,s256gat,s477gat);
  and x253(s1302gat,s256gat,s494gat);
  and x254(s1305gat,s256gat,s511gat);
  and x255(s1308gat,s256gat,s528gat);
  not x256(s1311gat,s591gat);
  not x257(s1315gat,s639gat);
  not x258(s1319gat,s687gat);
  not x259(s1323gat,s735gat);
  not x260(s1327gat,s783gat);
  not x261(s1331gat,s831gat);
  not x262(s1335gat,s879gat);
  not x263(s1339gat,s927gat);
  not x264(s1343gat,s975gat);
  not x265(s1347gat,s1023gat);
  not x266(s1351gat,s1071gat);
  not x267(s1355gat,s1119gat);
  not x268(s1359gat,s1167gat);
  not x269(s1363gat,s1215gat);
  not x270(s1367gat,s1263gat);
  nor x271(s1371gat,s591gat,s1311gat);
  not x272(s1372gat,s1311gat);
  nor x273(s1373gat,s639gat,s1315gat);
  not x274(s1374gat,s1315gat);
  nor x275(s1375gat,s687gat,s1319gat);
  not x276(s1376gat,s1319gat);
  nor x277(s1377gat,s735gat,s1323gat);
  not x278(s1378gat,s1323gat);
  nor x279(s1379gat,s783gat,s1327gat);
  not x280(s1380gat,s1327gat);
  nor x281(s1381gat,s831gat,s1331gat);
  not x282(s1382gat,s1331gat);
  nor x283(s1383gat,s879gat,s1335gat);
  not x284(s1384gat,s1335gat);
  nor x285(s1385gat,s927gat,s1339gat);
  not x286(s1386gat,s1339gat);
  nor x287(s1387gat,s975gat,s1343gat);
  not x288(s1388gat,s1343gat);
  nor x289(s1389gat,s1023gat,s1347gat);
  not x290(s1390gat,s1347gat);
  nor x291(s1391gat,s1071gat,s1351gat);
  not x292(s1392gat,s1351gat);
  nor x293(s1393gat,s1119gat,s1355gat);
  not x294(s1394gat,s1355gat);
  nor x295(s1395gat,s1167gat,s1359gat);
  not x296(s1396gat,s1359gat);
  nor x297(s1397gat,s1215gat,s1363gat);
  not x298(s1398gat,s1363gat);
  nor x299(s1399gat,s1263gat,s1367gat);
  not x300(s1400gat,s1367gat);
  nor x301(s1401gat,s1371gat,s1372gat);
  nor x302(s1404gat,s1373gat,s1374gat);
  nor x303(s1407gat,s1375gat,s1376gat);
  nor x304(s1410gat,s1377gat,s1378gat);
  nor x305(s1413gat,s1379gat,s1380gat);
  nor x306(s1416gat,s1381gat,s1382gat);
  nor x307(s1419gat,s1383gat,s1384gat);
  nor x308(s1422gat,s1385gat,s1386gat);
  nor x309(s1425gat,s1387gat,s1388gat);
  nor x310(s1428gat,s1389gat,s1390gat);
  nor x311(s1431gat,s1391gat,s1392gat);
  nor x312(s1434gat,s1393gat,s1394gat);
  nor x313(s1437gat,s1395gat,s1396gat);
  nor x314(s1440gat,s1397gat,s1398gat);
  nor x315(s1443gat,s1399gat,s1400gat);
  nor x316(s1446gat,s1401gat,s546gat);
  nor x317(s1450gat,s1404gat,s594gat);
  nor x318(s1454gat,s1407gat,s642gat);
  nor x319(s1458gat,s1410gat,s690gat);
  nor x320(s1462gat,s1413gat,s738gat);
  nor x321(s1466gat,s1416gat,s786gat);
  nor x322(s1470gat,s1419gat,s834gat);
  nor x323(s1474gat,s1422gat,s882gat);
  nor x324(s1478gat,s1425gat,s930gat);
  nor x325(s1482gat,s1428gat,s978gat);
  nor x326(s1486gat,s1431gat,s1026gat);
  nor x327(s1490gat,s1434gat,s1074gat);
  nor x328(s1494gat,s1437gat,s1122gat);
  nor x329(s1498gat,s1440gat,s1170gat);
  nor x330(s1502gat,s1443gat,s1218gat);
  nor x331(s1506gat,s1401gat,s1446gat);
  nor x332(s1507gat,s1446gat,s546gat);
  nor x333(s1508gat,s1311gat,s1446gat);
  nor x334(s1511gat,s1404gat,s1450gat);
  nor x335(s1512gat,s1450gat,s594gat);
  nor x336(s1513gat,s1315gat,s1450gat);
  nor x337(s1516gat,s1407gat,s1454gat);
  nor x338(s1517gat,s1454gat,s642gat);
  nor x339(s1518gat,s1319gat,s1454gat);
  nor x340(s1521gat,s1410gat,s1458gat);
  nor x341(s1522gat,s1458gat,s690gat);
  nor x342(s1523gat,s1323gat,s1458gat);
  nor x343(s1526gat,s1413gat,s1462gat);
  nor x344(s1527gat,s1462gat,s738gat);
  nor x345(s1528gat,s1327gat,s1462gat);
  nor x346(s1531gat,s1416gat,s1466gat);
  nor x347(s1532gat,s1466gat,s786gat);
  nor x348(s1533gat,s1331gat,s1466gat);
  nor x349(s1536gat,s1419gat,s1470gat);
  nor x350(s1537gat,s1470gat,s834gat);
  nor x351(s1538gat,s1335gat,s1470gat);
  nor x352(s1541gat,s1422gat,s1474gat);
  nor x353(s1542gat,s1474gat,s882gat);
  nor x354(s1543gat,s1339gat,s1474gat);
  nor x355(s1546gat,s1425gat,s1478gat);
  nor x356(s1547gat,s1478gat,s930gat);
  nor x357(s1548gat,s1343gat,s1478gat);
  nor x358(s1551gat,s1428gat,s1482gat);
  nor x359(s1552gat,s1482gat,s978gat);
  nor x360(s1553gat,s1347gat,s1482gat);
  nor x361(s1556gat,s1431gat,s1486gat);
  nor x362(s1557gat,s1486gat,s1026gat);
  nor x363(s1558gat,s1351gat,s1486gat);
  nor x364(s1561gat,s1434gat,s1490gat);
  nor x365(s1562gat,s1490gat,s1074gat);
  nor x366(s1563gat,s1355gat,s1490gat);
  nor x367(s1566gat,s1437gat,s1494gat);
  nor x368(s1567gat,s1494gat,s1122gat);
  nor x369(s1568gat,s1359gat,s1494gat);
  nor x370(s1571gat,s1440gat,s1498gat);
  nor x371(s1572gat,s1498gat,s1170gat);
  nor x372(s1573gat,s1363gat,s1498gat);
  nor x373(s1576gat,s1443gat,s1502gat);
  nor x374(s1577gat,s1502gat,s1218gat);
  nor x375(s1578gat,s1367gat,s1502gat);
  nor x376(s1581gat,s1506gat,s1507gat);
  nor x377(s1582gat,s1511gat,s1512gat);
  nor x378(s1585gat,s1516gat,s1517gat);
  nor x379(s1588gat,s1521gat,s1522gat);
  nor x380(s1591gat,s1526gat,s1527gat);
  nor x381(s1594gat,s1531gat,s1532gat);
  nor x382(s1597gat,s1536gat,s1537gat);
  nor x383(s1600gat,s1541gat,s1542gat);
  nor x384(s1603gat,s1546gat,s1547gat);
  nor x385(s1606gat,s1551gat,s1552gat);
  nor x386(s1609gat,s1556gat,s1557gat);
  nor x387(s1612gat,s1561gat,s1562gat);
  nor x388(s1615gat,s1566gat,s1567gat);
  nor x389(s1618gat,s1571gat,s1572gat);
  nor x390(s1621gat,s1576gat,s1577gat);
  nor x391(s1624gat,s1266gat,s1578gat);
  nor x392(s1628gat,s1582gat,s1508gat);
  nor x393(s1632gat,s1585gat,s1513gat);
  nor x394(s1636gat,s1588gat,s1518gat);
  nor x395(s1640gat,s1591gat,s1523gat);
  nor x396(s1644gat,s1594gat,s1528gat);
  nor x397(s1648gat,s1597gat,s1533gat);
  nor x398(s1652gat,s1600gat,s1538gat);
  nor x399(s1656gat,s1603gat,s1543gat);
  nor x400(s1660gat,s1606gat,s1548gat);
  nor x401(s1664gat,s1609gat,s1553gat);
  nor x402(s1668gat,s1612gat,s1558gat);
  nor x403(s1672gat,s1615gat,s1563gat);
  nor x404(s1676gat,s1618gat,s1568gat);
  nor x405(s1680gat,s1621gat,s1573gat);
  nor x406(s1684gat,s1266gat,s1624gat);
  nor x407(s1685gat,s1624gat,s1578gat);
  nor x408(s1686gat,s1582gat,s1628gat);
  nor x409(s1687gat,s1628gat,s1508gat);
  nor x410(s1688gat,s1585gat,s1632gat);
  nor x411(s1689gat,s1632gat,s1513gat);
  nor x412(s1690gat,s1588gat,s1636gat);
  nor x413(s1691gat,s1636gat,s1518gat);
  nor x414(s1692gat,s1591gat,s1640gat);
  nor x415(s1693gat,s1640gat,s1523gat);
  nor x416(s1694gat,s1594gat,s1644gat);
  nor x417(s1695gat,s1644gat,s1528gat);
  nor x418(s1696gat,s1597gat,s1648gat);
  nor x419(s1697gat,s1648gat,s1533gat);
  nor x420(s1698gat,s1600gat,s1652gat);
  nor x421(s1699gat,s1652gat,s1538gat);
  nor x422(s1700gat,s1603gat,s1656gat);
  nor x423(s1701gat,s1656gat,s1543gat);
  nor x424(s1702gat,s1606gat,s1660gat);
  nor x425(s1703gat,s1660gat,s1548gat);
  nor x426(s1704gat,s1609gat,s1664gat);
  nor x427(s1705gat,s1664gat,s1553gat);
  nor x428(s1706gat,s1612gat,s1668gat);
  nor x429(s1707gat,s1668gat,s1558gat);
  nor x430(s1708gat,s1615gat,s1672gat);
  nor x431(s1709gat,s1672gat,s1563gat);
  nor x432(s1710gat,s1618gat,s1676gat);
  nor x433(s1711gat,s1676gat,s1568gat);
  nor x434(s1712gat,s1621gat,s1680gat);
  nor x435(s1713gat,s1680gat,s1573gat);
  nor x436(s1714gat,s1684gat,s1685gat);
  nor x437(s1717gat,s1686gat,s1687gat);
  nor x438(s1720gat,s1688gat,s1689gat);
  nor x439(s1723gat,s1690gat,s1691gat);
  nor x440(s1726gat,s1692gat,s1693gat);
  nor x441(s1729gat,s1694gat,s1695gat);
  nor x442(s1732gat,s1696gat,s1697gat);
  nor x443(s1735gat,s1698gat,s1699gat);
  nor x444(s1738gat,s1700gat,s1701gat);
  nor x445(s1741gat,s1702gat,s1703gat);
  nor x446(s1744gat,s1704gat,s1705gat);
  nor x447(s1747gat,s1706gat,s1707gat);
  nor x448(s1750gat,s1708gat,s1709gat);
  nor x449(s1753gat,s1710gat,s1711gat);
  nor x450(s1756gat,s1712gat,s1713gat);
  nor x451(s1759gat,s1714gat,s1221gat);
  nor x452(s1763gat,s1717gat,s549gat);
  nor x453(s1767gat,s1720gat,s597gat);
  nor x454(s1771gat,s1723gat,s645gat);
  nor x455(s1775gat,s1726gat,s693gat);
  nor x456(s1779gat,s1729gat,s741gat);
  nor x457(s1783gat,s1732gat,s789gat);
  nor x458(s1787gat,s1735gat,s837gat);
  nor x459(s1791gat,s1738gat,s885gat);
  nor x460(s1795gat,s1741gat,s933gat);
  nor x461(s1799gat,s1744gat,s981gat);
  nor x462(s1803gat,s1747gat,s1029gat);
  nor x463(s1807gat,s1750gat,s1077gat);
  nor x464(s1811gat,s1753gat,s1125gat);
  nor x465(s1815gat,s1756gat,s1173gat);
  nor x466(s1819gat,s1714gat,s1759gat);
  nor x467(s1820gat,s1759gat,s1221gat);
  nor x468(s1821gat,s1624gat,s1759gat);
  nor x469(s1824gat,s1717gat,s1763gat);
  nor x470(s1825gat,s1763gat,s549gat);
  nor x471(s1826gat,s1628gat,s1763gat);
  nor x472(s1829gat,s1720gat,s1767gat);
  nor x473(s1830gat,s1767gat,s597gat);
  nor x474(s1831gat,s1632gat,s1767gat);
  nor x475(s1834gat,s1723gat,s1771gat);
  nor x476(s1835gat,s1771gat,s645gat);
  nor x477(s1836gat,s1636gat,s1771gat);
  nor x478(s1839gat,s1726gat,s1775gat);
  nor x479(s1840gat,s1775gat,s693gat);
  nor x480(s1841gat,s1640gat,s1775gat);
  nor x481(s1844gat,s1729gat,s1779gat);
  nor x482(s1845gat,s1779gat,s741gat);
  nor x483(s1846gat,s1644gat,s1779gat);
  nor x484(s1849gat,s1732gat,s1783gat);
  nor x485(s1850gat,s1783gat,s789gat);
  nor x486(s1851gat,s1648gat,s1783gat);
  nor x487(s1854gat,s1735gat,s1787gat);
  nor x488(s1855gat,s1787gat,s837gat);
  nor x489(s1856gat,s1652gat,s1787gat);
  nor x490(s1859gat,s1738gat,s1791gat);
  nor x491(s1860gat,s1791gat,s885gat);
  nor x492(s1861gat,s1656gat,s1791gat);
  nor x493(s1864gat,s1741gat,s1795gat);
  nor x494(s1865gat,s1795gat,s933gat);
  nor x495(s1866gat,s1660gat,s1795gat);
  nor x496(s1869gat,s1744gat,s1799gat);
  nor x497(s1870gat,s1799gat,s981gat);
  nor x498(s1871gat,s1664gat,s1799gat);
  nor x499(s1874gat,s1747gat,s1803gat);
  nor x500(s1875gat,s1803gat,s1029gat);
  nor x501(s1876gat,s1668gat,s1803gat);
  nor x502(s1879gat,s1750gat,s1807gat);
  nor x503(s1880gat,s1807gat,s1077gat);
  nor x504(s1881gat,s1672gat,s1807gat);
  nor x505(s1884gat,s1753gat,s1811gat);
  nor x506(s1885gat,s1811gat,s1125gat);
  nor x507(s1886gat,s1676gat,s1811gat);
  nor x508(s1889gat,s1756gat,s1815gat);
  nor x509(s1890gat,s1815gat,s1173gat);
  nor x510(s1891gat,s1680gat,s1815gat);
  nor x511(s1894gat,s1819gat,s1820gat);
  nor x512(s1897gat,s1269gat,s1821gat);
  nor x513(s1901gat,s1824gat,s1825gat);
  nor x514(s1902gat,s1829gat,s1830gat);
  nor x515(s1905gat,s1834gat,s1835gat);
  nor x516(s1908gat,s1839gat,s1840gat);
  nor x517(s1911gat,s1844gat,s1845gat);
  nor x518(s1914gat,s1849gat,s1850gat);
  nor x519(s1917gat,s1854gat,s1855gat);
  nor x520(s1920gat,s1859gat,s1860gat);
  nor x521(s1923gat,s1864gat,s1865gat);
  nor x522(s1926gat,s1869gat,s1870gat);
  nor x523(s1929gat,s1874gat,s1875gat);
  nor x524(s1932gat,s1879gat,s1880gat);
  nor x525(s1935gat,s1884gat,s1885gat);
  nor x526(s1938gat,s1889gat,s1890gat);
  nor x527(s1941gat,s1894gat,s1891gat);
  nor x528(s1945gat,s1269gat,s1897gat);
  nor x529(s1946gat,s1897gat,s1821gat);
  nor x530(s1947gat,s1902gat,s1826gat);
  nor x531(s1951gat,s1905gat,s1831gat);
  nor x532(s1955gat,s1908gat,s1836gat);
  nor x533(s1959gat,s1911gat,s1841gat);
  nor x534(s1963gat,s1914gat,s1846gat);
  nor x535(s1967gat,s1917gat,s1851gat);
  nor x536(s1971gat,s1920gat,s1856gat);
  nor x537(s1975gat,s1923gat,s1861gat);
  nor x538(s1979gat,s1926gat,s1866gat);
  nor x539(s1983gat,s1929gat,s1871gat);
  nor x540(s1987gat,s1932gat,s1876gat);
  nor x541(s1991gat,s1935gat,s1881gat);
  nor x542(s1995gat,s1938gat,s1886gat);
  nor x543(s1999gat,s1894gat,s1941gat);
  nor x544(s2000gat,s1941gat,s1891gat);
  nor x545(s2001gat,s1945gat,s1946gat);
  nor x546(s2004gat,s1902gat,s1947gat);
  nor x547(s2005gat,s1947gat,s1826gat);
  nor x548(s2006gat,s1905gat,s1951gat);
  nor x549(s2007gat,s1951gat,s1831gat);
  nor x550(s2008gat,s1908gat,s1955gat);
  nor x551(s2009gat,s1955gat,s1836gat);
  nor x552(s2010gat,s1911gat,s1959gat);
  nor x553(s2011gat,s1959gat,s1841gat);
  nor x554(s2012gat,s1914gat,s1963gat);
  nor x555(s2013gat,s1963gat,s1846gat);
  nor x556(s2014gat,s1917gat,s1967gat);
  nor x557(s2015gat,s1967gat,s1851gat);
  nor x558(s2016gat,s1920gat,s1971gat);
  nor x559(s2017gat,s1971gat,s1856gat);
  nor x560(s2018gat,s1923gat,s1975gat);
  nor x561(s2019gat,s1975gat,s1861gat);
  nor x562(s2020gat,s1926gat,s1979gat);
  nor x563(s2021gat,s1979gat,s1866gat);
  nor x564(s2022gat,s1929gat,s1983gat);
  nor x565(s2023gat,s1983gat,s1871gat);
  nor x566(s2024gat,s1932gat,s1987gat);
  nor x567(s2025gat,s1987gat,s1876gat);
  nor x568(s2026gat,s1935gat,s1991gat);
  nor x569(s2027gat,s1991gat,s1881gat);
  nor x570(s2028gat,s1938gat,s1995gat);
  nor x571(s2029gat,s1995gat,s1886gat);
  nor x572(s2030gat,s1999gat,s2000gat);
  nor x573(s2033gat,s2001gat,s1224gat);
  nor x574(s2037gat,s2004gat,s2005gat);
  nor x575(s2040gat,s2006gat,s2007gat);
  nor x576(s2043gat,s2008gat,s2009gat);
  nor x577(s2046gat,s2010gat,s2011gat);
  nor x578(s2049gat,s2012gat,s2013gat);
  nor x579(s2052gat,s2014gat,s2015gat);
  nor x580(s2055gat,s2016gat,s2017gat);
  nor x581(s2058gat,s2018gat,s2019gat);
  nor x582(s2061gat,s2020gat,s2021gat);
  nor x583(s2064gat,s2022gat,s2023gat);
  nor x584(s2067gat,s2024gat,s2025gat);
  nor x585(s2070gat,s2026gat,s2027gat);
  nor x586(s2073gat,s2028gat,s2029gat);
  nor x587(s2076gat,s2030gat,s1176gat);
  nor x588(s2080gat,s2001gat,s2033gat);
  nor x589(s2081gat,s2033gat,s1224gat);
  nor x590(s2082gat,s1897gat,s2033gat);
  nor x591(s2085gat,s2037gat,s552gat);
  nor x592(s2089gat,s2040gat,s600gat);
  nor x593(s2093gat,s2043gat,s648gat);
  nor x594(s2097gat,s2046gat,s696gat);
  nor x595(s2101gat,s2049gat,s744gat);
  nor x596(s2105gat,s2052gat,s792gat);
  nor x597(s2109gat,s2055gat,s840gat);
  nor x598(s2113gat,s2058gat,s888gat);
  nor x599(s2117gat,s2061gat,s936gat);
  nor x600(s2121gat,s2064gat,s984gat);
  nor x601(s2125gat,s2067gat,s1032gat);
  nor x602(s2129gat,s2070gat,s1080gat);
  nor x603(s2133gat,s2073gat,s1128gat);
  nor x604(s2137gat,s2030gat,s2076gat);
  nor x605(s2138gat,s2076gat,s1176gat);
  nor x606(s2139gat,s1941gat,s2076gat);
  nor x607(s2142gat,s2080gat,s2081gat);
  nor x608(s2145gat,s1272gat,s2082gat);
  nor x609(s2149gat,s2037gat,s2085gat);
  nor x610(s2150gat,s2085gat,s552gat);
  nor x611(s2151gat,s1947gat,s2085gat);
  nor x612(s2154gat,s2040gat,s2089gat);
  nor x613(s2155gat,s2089gat,s600gat);
  nor x614(s2156gat,s1951gat,s2089gat);
  nor x615(s2159gat,s2043gat,s2093gat);
  nor x616(s2160gat,s2093gat,s648gat);
  nor x617(s2161gat,s1955gat,s2093gat);
  nor x618(s2164gat,s2046gat,s2097gat);
  nor x619(s2165gat,s2097gat,s696gat);
  nor x620(s2166gat,s1959gat,s2097gat);
  nor x621(s2169gat,s2049gat,s2101gat);
  nor x622(s2170gat,s2101gat,s744gat);
  nor x623(s2171gat,s1963gat,s2101gat);
  nor x624(s2174gat,s2052gat,s2105gat);
  nor x625(s2175gat,s2105gat,s792gat);
  nor x626(s2176gat,s1967gat,s2105gat);
  nor x627(s2179gat,s2055gat,s2109gat);
  nor x628(s2180gat,s2109gat,s840gat);
  nor x629(s2181gat,s1971gat,s2109gat);
  nor x630(s2184gat,s2058gat,s2113gat);
  nor x631(s2185gat,s2113gat,s888gat);
  nor x632(s2186gat,s1975gat,s2113gat);
  nor x633(s2189gat,s2061gat,s2117gat);
  nor x634(s2190gat,s2117gat,s936gat);
  nor x635(s2191gat,s1979gat,s2117gat);
  nor x636(s2194gat,s2064gat,s2121gat);
  nor x637(s2195gat,s2121gat,s984gat);
  nor x638(s2196gat,s1983gat,s2121gat);
  nor x639(s2199gat,s2067gat,s2125gat);
  nor x640(s2200gat,s2125gat,s1032gat);
  nor x641(s2201gat,s1987gat,s2125gat);
  nor x642(s2204gat,s2070gat,s2129gat);
  nor x643(s2205gat,s2129gat,s1080gat);
  nor x644(s2206gat,s1991gat,s2129gat);
  nor x645(s2209gat,s2073gat,s2133gat);
  nor x646(s2210gat,s2133gat,s1128gat);
  nor x647(s2211gat,s1995gat,s2133gat);
  nor x648(s2214gat,s2137gat,s2138gat);
  nor x649(s2217gat,s2142gat,s2139gat);
  nor x650(s2221gat,s1272gat,s2145gat);
  nor x651(s2222gat,s2145gat,s2082gat);
  nor x652(s2223gat,s2149gat,s2150gat);
  nor x653(s2224gat,s2154gat,s2155gat);
  nor x654(s2227gat,s2159gat,s2160gat);
  nor x655(s2230gat,s2164gat,s2165gat);
  nor x656(s2233gat,s2169gat,s2170gat);
  nor x657(s2236gat,s2174gat,s2175gat);
  nor x658(s2239gat,s2179gat,s2180gat);
  nor x659(s2242gat,s2184gat,s2185gat);
  nor x660(s2245gat,s2189gat,s2190gat);
  nor x661(s2248gat,s2194gat,s2195gat);
  nor x662(s2251gat,s2199gat,s2200gat);
  nor x663(s2254gat,s2204gat,s2205gat);
  nor x664(s2257gat,s2209gat,s2210gat);
  nor x665(s2260gat,s2214gat,s2211gat);
  nor x666(s2264gat,s2142gat,s2217gat);
  nor x667(s2265gat,s2217gat,s2139gat);
  nor x668(s2266gat,s2221gat,s2222gat);
  nor x669(s2269gat,s2224gat,s2151gat);
  nor x670(s2273gat,s2227gat,s2156gat);
  nor x671(s2277gat,s2230gat,s2161gat);
  nor x672(s2281gat,s2233gat,s2166gat);
  nor x673(s2285gat,s2236gat,s2171gat);
  nor x674(s2289gat,s2239gat,s2176gat);
  nor x675(s2293gat,s2242gat,s2181gat);
  nor x676(s2297gat,s2245gat,s2186gat);
  nor x677(s2301gat,s2248gat,s2191gat);
  nor x678(s2305gat,s2251gat,s2196gat);
  nor x679(s2309gat,s2254gat,s2201gat);
  nor x680(s2313gat,s2257gat,s2206gat);
  nor x681(s2317gat,s2214gat,s2260gat);
  nor x682(s2318gat,s2260gat,s2211gat);
  nor x683(s2319gat,s2264gat,s2265gat);
  nor x684(s2322gat,s2266gat,s1227gat);
  nor x685(s2326gat,s2224gat,s2269gat);
  nor x686(s2327gat,s2269gat,s2151gat);
  nor x687(s2328gat,s2227gat,s2273gat);
  nor x688(s2329gat,s2273gat,s2156gat);
  nor x689(s2330gat,s2230gat,s2277gat);
  nor x690(s2331gat,s2277gat,s2161gat);
  nor x691(s2332gat,s2233gat,s2281gat);
  nor x692(s2333gat,s2281gat,s2166gat);
  nor x693(s2334gat,s2236gat,s2285gat);
  nor x694(s2335gat,s2285gat,s2171gat);
  nor x695(s2336gat,s2239gat,s2289gat);
  nor x696(s2337gat,s2289gat,s2176gat);
  nor x697(s2338gat,s2242gat,s2293gat);
  nor x698(s2339gat,s2293gat,s2181gat);
  nor x699(s2340gat,s2245gat,s2297gat);
  nor x700(s2341gat,s2297gat,s2186gat);
  nor x701(s2342gat,s2248gat,s2301gat);
  nor x702(s2343gat,s2301gat,s2191gat);
  nor x703(s2344gat,s2251gat,s2305gat);
  nor x704(s2345gat,s2305gat,s2196gat);
  nor x705(s2346gat,s2254gat,s2309gat);
  nor x706(s2347gat,s2309gat,s2201gat);
  nor x707(s2348gat,s2257gat,s2313gat);
  nor x708(s2349gat,s2313gat,s2206gat);
  nor x709(s2350gat,s2317gat,s2318gat);
  nor x710(s2353gat,s2319gat,s1179gat);
  nor x711(s2357gat,s2266gat,s2322gat);
  nor x712(s2358gat,s2322gat,s1227gat);
  nor x713(s2359gat,s2145gat,s2322gat);
  nor x714(s2362gat,s2326gat,s2327gat);
  nor x715(s2365gat,s2328gat,s2329gat);
  nor x716(s2368gat,s2330gat,s2331gat);
  nor x717(s2371gat,s2332gat,s2333gat);
  nor x718(s2374gat,s2334gat,s2335gat);
  nor x719(s2377gat,s2336gat,s2337gat);
  nor x720(s2380gat,s2338gat,s2339gat);
  nor x721(s2383gat,s2340gat,s2341gat);
  nor x722(s2386gat,s2342gat,s2343gat);
  nor x723(s2389gat,s2344gat,s2345gat);
  nor x724(s2392gat,s2346gat,s2347gat);
  nor x725(s2395gat,s2348gat,s2349gat);
  nor x726(s2398gat,s2350gat,s1131gat);
  nor x727(s2402gat,s2319gat,s2353gat);
  nor x728(s2403gat,s2353gat,s1179gat);
  nor x729(s2404gat,s2217gat,s2353gat);
  nor x730(s2407gat,s2357gat,s2358gat);
  nor x731(s2410gat,s1275gat,s2359gat);
  nor x732(s2414gat,s2362gat,s555gat);
  nor x733(s2418gat,s2365gat,s603gat);
  nor x734(s2422gat,s2368gat,s651gat);
  nor x735(s2426gat,s2371gat,s699gat);
  nor x736(s2430gat,s2374gat,s747gat);
  nor x737(s2434gat,s2377gat,s795gat);
  nor x738(s2438gat,s2380gat,s843gat);
  nor x739(s2442gat,s2383gat,s891gat);
  nor x740(s2446gat,s2386gat,s939gat);
  nor x741(s2450gat,s2389gat,s987gat);
  nor x742(s2454gat,s2392gat,s1035gat);
  nor x743(s2458gat,s2395gat,s1083gat);
  nor x744(s2462gat,s2350gat,s2398gat);
  nor x745(s2463gat,s2398gat,s1131gat);
  nor x746(s2464gat,s2260gat,s2398gat);
  nor x747(s2467gat,s2402gat,s2403gat);
  nor x748(s2470gat,s2407gat,s2404gat);
  nor x749(s2474gat,s1275gat,s2410gat);
  nor x750(s2475gat,s2410gat,s2359gat);
  nor x751(s2476gat,s2362gat,s2414gat);
  nor x752(s2477gat,s2414gat,s555gat);
  nor x753(s2478gat,s2269gat,s2414gat);
  nor x754(s2481gat,s2365gat,s2418gat);
  nor x755(s2482gat,s2418gat,s603gat);
  nor x756(s2483gat,s2273gat,s2418gat);
  nor x757(s2486gat,s2368gat,s2422gat);
  nor x758(s2487gat,s2422gat,s651gat);
  nor x759(s2488gat,s2277gat,s2422gat);
  nor x760(s2491gat,s2371gat,s2426gat);
  nor x761(s2492gat,s2426gat,s699gat);
  nor x762(s2493gat,s2281gat,s2426gat);
  nor x763(s2496gat,s2374gat,s2430gat);
  nor x764(s2497gat,s2430gat,s747gat);
  nor x765(s2498gat,s2285gat,s2430gat);
  nor x766(s2501gat,s2377gat,s2434gat);
  nor x767(s2502gat,s2434gat,s795gat);
  nor x768(s2503gat,s2289gat,s2434gat);
  nor x769(s2506gat,s2380gat,s2438gat);
  nor x770(s2507gat,s2438gat,s843gat);
  nor x771(s2508gat,s2293gat,s2438gat);
  nor x772(s2511gat,s2383gat,s2442gat);
  nor x773(s2512gat,s2442gat,s891gat);
  nor x774(s2513gat,s2297gat,s2442gat);
  nor x775(s2516gat,s2386gat,s2446gat);
  nor x776(s2517gat,s2446gat,s939gat);
  nor x777(s2518gat,s2301gat,s2446gat);
  nor x778(s2521gat,s2389gat,s2450gat);
  nor x779(s2522gat,s2450gat,s987gat);
  nor x780(s2523gat,s2305gat,s2450gat);
  nor x781(s2526gat,s2392gat,s2454gat);
  nor x782(s2527gat,s2454gat,s1035gat);
  nor x783(s2528gat,s2309gat,s2454gat);
  nor x784(s2531gat,s2395gat,s2458gat);
  nor x785(s2532gat,s2458gat,s1083gat);
  nor x786(s2533gat,s2313gat,s2458gat);
  nor x787(s2536gat,s2462gat,s2463gat);
  nor x788(s2539gat,s2467gat,s2464gat);
  nor x789(s2543gat,s2407gat,s2470gat);
  nor x790(s2544gat,s2470gat,s2404gat);
  nor x791(s2545gat,s2474gat,s2475gat);
  nor x792(s2548gat,s2476gat,s2477gat);
  nor x793(s2549gat,s2481gat,s2482gat);
  nor x794(s2552gat,s2486gat,s2487gat);
  nor x795(s2555gat,s2491gat,s2492gat);
  nor x796(s2558gat,s2496gat,s2497gat);
  nor x797(s2561gat,s2501gat,s2502gat);
  nor x798(s2564gat,s2506gat,s2507gat);
  nor x799(s2567gat,s2511gat,s2512gat);
  nor x800(s2570gat,s2516gat,s2517gat);
  nor x801(s2573gat,s2521gat,s2522gat);
  nor x802(s2576gat,s2526gat,s2527gat);
  nor x803(s2579gat,s2531gat,s2532gat);
  nor x804(s2582gat,s2536gat,s2533gat);
  nor x805(s2586gat,s2467gat,s2539gat);
  nor x806(s2587gat,s2539gat,s2464gat);
  nor x807(s2588gat,s2543gat,s2544gat);
  nor x808(s2591gat,s2545gat,s1230gat);
  nor x809(s2595gat,s2549gat,s2478gat);
  nor x810(s2599gat,s2552gat,s2483gat);
  nor x811(s2603gat,s2555gat,s2488gat);
  nor x812(s2607gat,s2558gat,s2493gat);
  nor x813(s2611gat,s2561gat,s2498gat);
  nor x814(s2615gat,s2564gat,s2503gat);
  nor x815(s2619gat,s2567gat,s2508gat);
  nor x816(s2623gat,s2570gat,s2513gat);
  nor x817(s2627gat,s2573gat,s2518gat);
  nor x818(s2631gat,s2576gat,s2523gat);
  nor x819(s2635gat,s2579gat,s2528gat);
  nor x820(s2639gat,s2536gat,s2582gat);
  nor x821(s2640gat,s2582gat,s2533gat);
  nor x822(s2641gat,s2586gat,s2587gat);
  nor x823(s2644gat,s2588gat,s1182gat);
  nor x824(s2648gat,s2545gat,s2591gat);
  nor x825(s2649gat,s2591gat,s1230gat);
  nor x826(s2650gat,s2410gat,s2591gat);
  nor x827(s2653gat,s2549gat,s2595gat);
  nor x828(s2654gat,s2595gat,s2478gat);
  nor x829(s2655gat,s2552gat,s2599gat);
  nor x830(s2656gat,s2599gat,s2483gat);
  nor x831(s2657gat,s2555gat,s2603gat);
  nor x832(s2658gat,s2603gat,s2488gat);
  nor x833(s2659gat,s2558gat,s2607gat);
  nor x834(s2660gat,s2607gat,s2493gat);
  nor x835(s2661gat,s2561gat,s2611gat);
  nor x836(s2662gat,s2611gat,s2498gat);
  nor x837(s2663gat,s2564gat,s2615gat);
  nor x838(s2664gat,s2615gat,s2503gat);
  nor x839(s2665gat,s2567gat,s2619gat);
  nor x840(s2666gat,s2619gat,s2508gat);
  nor x841(s2667gat,s2570gat,s2623gat);
  nor x842(s2668gat,s2623gat,s2513gat);
  nor x843(s2669gat,s2573gat,s2627gat);
  nor x844(s2670gat,s2627gat,s2518gat);
  nor x845(s2671gat,s2576gat,s2631gat);
  nor x846(s2672gat,s2631gat,s2523gat);
  nor x847(s2673gat,s2579gat,s2635gat);
  nor x848(s2674gat,s2635gat,s2528gat);
  nor x849(s2675gat,s2639gat,s2640gat);
  nor x850(s2678gat,s2641gat,s1134gat);
  nor x851(s2682gat,s2588gat,s2644gat);
  nor x852(s2683gat,s2644gat,s1182gat);
  nor x853(s2684gat,s2470gat,s2644gat);
  nor x854(s2687gat,s2648gat,s2649gat);
  nor x855(s2690gat,s1278gat,s2650gat);
  nor x856(s2694gat,s2653gat,s2654gat);
  nor x857(s2697gat,s2655gat,s2656gat);
  nor x858(s2700gat,s2657gat,s2658gat);
  nor x859(s2703gat,s2659gat,s2660gat);
  nor x860(s2706gat,s2661gat,s2662gat);
  nor x861(s2709gat,s2663gat,s2664gat);
  nor x862(s2712gat,s2665gat,s2666gat);
  nor x863(s2715gat,s2667gat,s2668gat);
  nor x864(s2718gat,s2669gat,s2670gat);
  nor x865(s2721gat,s2671gat,s2672gat);
  nor x866(s2724gat,s2673gat,s2674gat);
  nor x867(s2727gat,s2675gat,s1086gat);
  nor x868(s2731gat,s2641gat,s2678gat);
  nor x869(s2732gat,s2678gat,s1134gat);
  nor x870(s2733gat,s2539gat,s2678gat);
  nor x871(s2736gat,s2682gat,s2683gat);
  nor x872(s2739gat,s2687gat,s2684gat);
  nor x873(s2743gat,s1278gat,s2690gat);
  nor x874(s2744gat,s2690gat,s2650gat);
  nor x875(s2745gat,s2694gat,s558gat);
  nor x876(s2749gat,s2697gat,s606gat);
  nor x877(s2753gat,s2700gat,s654gat);
  nor x878(s2757gat,s2703gat,s702gat);
  nor x879(s2761gat,s2706gat,s750gat);
  nor x880(s2765gat,s2709gat,s798gat);
  nor x881(s2769gat,s2712gat,s846gat);
  nor x882(s2773gat,s2715gat,s894gat);
  nor x883(s2777gat,s2718gat,s942gat);
  nor x884(s2781gat,s2721gat,s990gat);
  nor x885(s2785gat,s2724gat,s1038gat);
  nor x886(s2789gat,s2675gat,s2727gat);
  nor x887(s2790gat,s2727gat,s1086gat);
  nor x888(s2791gat,s2582gat,s2727gat);
  nor x889(s2794gat,s2731gat,s2732gat);
  nor x890(s2797gat,s2736gat,s2733gat);
  nor x891(s2801gat,s2687gat,s2739gat);
  nor x892(s2802gat,s2739gat,s2684gat);
  nor x893(s2803gat,s2743gat,s2744gat);
  nor x894(s2806gat,s2694gat,s2745gat);
  nor x895(s2807gat,s2745gat,s558gat);
  nor x896(s2808gat,s2595gat,s2745gat);
  nor x897(s2811gat,s2697gat,s2749gat);
  nor x898(s2812gat,s2749gat,s606gat);
  nor x899(s2813gat,s2599gat,s2749gat);
  nor x900(s2816gat,s2700gat,s2753gat);
  nor x901(s2817gat,s2753gat,s654gat);
  nor x902(s2818gat,s2603gat,s2753gat);
  nor x903(s2821gat,s2703gat,s2757gat);
  nor x904(s2822gat,s2757gat,s702gat);
  nor x905(s2823gat,s2607gat,s2757gat);
  nor x906(s2826gat,s2706gat,s2761gat);
  nor x907(s2827gat,s2761gat,s750gat);
  nor x908(s2828gat,s2611gat,s2761gat);
  nor x909(s2831gat,s2709gat,s2765gat);
  nor x910(s2832gat,s2765gat,s798gat);
  nor x911(s2833gat,s2615gat,s2765gat);
  nor x912(s2836gat,s2712gat,s2769gat);
  nor x913(s2837gat,s2769gat,s846gat);
  nor x914(s2838gat,s2619gat,s2769gat);
  nor x915(s2841gat,s2715gat,s2773gat);
  nor x916(s2842gat,s2773gat,s894gat);
  nor x917(s2843gat,s2623gat,s2773gat);
  nor x918(s2846gat,s2718gat,s2777gat);
  nor x919(s2847gat,s2777gat,s942gat);
  nor x920(s2848gat,s2627gat,s2777gat);
  nor x921(s2851gat,s2721gat,s2781gat);
  nor x922(s2852gat,s2781gat,s990gat);
  nor x923(s2853gat,s2631gat,s2781gat);
  nor x924(s2856gat,s2724gat,s2785gat);
  nor x925(s2857gat,s2785gat,s1038gat);
  nor x926(s2858gat,s2635gat,s2785gat);
  nor x927(s2861gat,s2789gat,s2790gat);
  nor x928(s2864gat,s2794gat,s2791gat);
  nor x929(s2868gat,s2736gat,s2797gat);
  nor x930(s2869gat,s2797gat,s2733gat);
  nor x931(s2870gat,s2801gat,s2802gat);
  nor x932(s2873gat,s2803gat,s1233gat);
  nor x933(s2877gat,s2806gat,s2807gat);
  nor x934(s2878gat,s2811gat,s2812gat);
  nor x935(s2881gat,s2816gat,s2817gat);
  nor x936(s2884gat,s2821gat,s2822gat);
  nor x937(s2887gat,s2826gat,s2827gat);
  nor x938(s2890gat,s2831gat,s2832gat);
  nor x939(s2893gat,s2836gat,s2837gat);
  nor x940(s2896gat,s2841gat,s2842gat);
  nor x941(s2899gat,s2846gat,s2847gat);
  nor x942(s2902gat,s2851gat,s2852gat);
  nor x943(s2905gat,s2856gat,s2857gat);
  nor x944(s2908gat,s2861gat,s2858gat);
  nor x945(s2912gat,s2794gat,s2864gat);
  nor x946(s2913gat,s2864gat,s2791gat);
  nor x947(s2914gat,s2868gat,s2869gat);
  nor x948(s2917gat,s2870gat,s1185gat);
  nor x949(s2921gat,s2803gat,s2873gat);
  nor x950(s2922gat,s2873gat,s1233gat);
  nor x951(s2923gat,s2690gat,s2873gat);
  nor x952(s2926gat,s2878gat,s2808gat);
  nor x953(s2930gat,s2881gat,s2813gat);
  nor x954(s2934gat,s2884gat,s2818gat);
  nor x955(s2938gat,s2887gat,s2823gat);
  nor x956(s2942gat,s2890gat,s2828gat);
  nor x957(s2946gat,s2893gat,s2833gat);
  nor x958(s2950gat,s2896gat,s2838gat);
  nor x959(s2954gat,s2899gat,s2843gat);
  nor x960(s2958gat,s2902gat,s2848gat);
  nor x961(s2962gat,s2905gat,s2853gat);
  nor x962(s2966gat,s2861gat,s2908gat);
  nor x963(s2967gat,s2908gat,s2858gat);
  nor x964(s2968gat,s2912gat,s2913gat);
  nor x965(s2971gat,s2914gat,s1137gat);
  nor x966(s2975gat,s2870gat,s2917gat);
  nor x967(s2976gat,s2917gat,s1185gat);
  nor x968(s2977gat,s2739gat,s2917gat);
  nor x969(s2980gat,s2921gat,s2922gat);
  nor x970(s2983gat,s1281gat,s2923gat);
  nor x971(s2987gat,s2878gat,s2926gat);
  nor x972(s2988gat,s2926gat,s2808gat);
  nor x973(s2989gat,s2881gat,s2930gat);
  nor x974(s2990gat,s2930gat,s2813gat);
  nor x975(s2991gat,s2884gat,s2934gat);
  nor x976(s2992gat,s2934gat,s2818gat);
  nor x977(s2993gat,s2887gat,s2938gat);
  nor x978(s2994gat,s2938gat,s2823gat);
  nor x979(s2995gat,s2890gat,s2942gat);
  nor x980(s2996gat,s2942gat,s2828gat);
  nor x981(s2997gat,s2893gat,s2946gat);
  nor x982(s2998gat,s2946gat,s2833gat);
  nor x983(s2999gat,s2896gat,s2950gat);
  nor x984(s3000gat,s2950gat,s2838gat);
  nor x985(s3001gat,s2899gat,s2954gat);
  nor x986(s3002gat,s2954gat,s2843gat);
  nor x987(s3003gat,s2902gat,s2958gat);
  nor x988(s3004gat,s2958gat,s2848gat);
  nor x989(s3005gat,s2905gat,s2962gat);
  nor x990(s3006gat,s2962gat,s2853gat);
  nor x991(s3007gat,s2966gat,s2967gat);
  nor x992(s3010gat,s2968gat,s1089gat);
  nor x993(s3014gat,s2914gat,s2971gat);
  nor x994(s3015gat,s2971gat,s1137gat);
  nor x995(s3016gat,s2797gat,s2971gat);
  nor x996(s3019gat,s2975gat,s2976gat);
  nor x997(s3022gat,s2980gat,s2977gat);
  nor x998(s3026gat,s1281gat,s2983gat);
  nor x999(s3027gat,s2983gat,s2923gat);
  nor x1000(s3028gat,s2987gat,s2988gat);
  nor x1001(s3031gat,s2989gat,s2990gat);
  nor x1002(s3034gat,s2991gat,s2992gat);
  nor x1003(s3037gat,s2993gat,s2994gat);
  nor x1004(s3040gat,s2995gat,s2996gat);
  nor x1005(s3043gat,s2997gat,s2998gat);
  nor x1006(s3046gat,s2999gat,s3000gat);
  nor x1007(s3049gat,s3001gat,s3002gat);
  nor x1008(s3052gat,s3003gat,s3004gat);
  nor x1009(s3055gat,s3005gat,s3006gat);
  nor x1010(s3058gat,s3007gat,s1041gat);
  nor x1011(s3062gat,s2968gat,s3010gat);
  nor x1012(s3063gat,s3010gat,s1089gat);
  nor x1013(s3064gat,s2864gat,s3010gat);
  nor x1014(s3067gat,s3014gat,s3015gat);
  nor x1015(s3070gat,s3019gat,s3016gat);
  nor x1016(s3074gat,s2980gat,s3022gat);
  nor x1017(s3075gat,s3022gat,s2977gat);
  nor x1018(s3076gat,s3026gat,s3027gat);
  nor x1019(s3079gat,s3028gat,s561gat);
  nor x1020(s3083gat,s3031gat,s609gat);
  nor x1021(s3087gat,s3034gat,s657gat);
  nor x1022(s3091gat,s3037gat,s705gat);
  nor x1023(s3095gat,s3040gat,s753gat);
  nor x1024(s3099gat,s3043gat,s801gat);
  nor x1025(s3103gat,s3046gat,s849gat);
  nor x1026(s3107gat,s3049gat,s897gat);
  nor x1027(s3111gat,s3052gat,s945gat);
  nor x1028(s3115gat,s3055gat,s993gat);
  nor x1029(s3119gat,s3007gat,s3058gat);
  nor x1030(s3120gat,s3058gat,s1041gat);
  nor x1031(s3121gat,s2908gat,s3058gat);
  nor x1032(s3124gat,s3062gat,s3063gat);
  nor x1033(s3127gat,s3067gat,s3064gat);
  nor x1034(s3131gat,s3019gat,s3070gat);
  nor x1035(s3132gat,s3070gat,s3016gat);
  nor x1036(s3133gat,s3074gat,s3075gat);
  nor x1037(s3136gat,s3076gat,s1236gat);
  nor x1038(s3140gat,s3028gat,s3079gat);
  nor x1039(s3141gat,s3079gat,s561gat);
  nor x1040(s3142gat,s2926gat,s3079gat);
  nor x1041(s3145gat,s3031gat,s3083gat);
  nor x1042(s3146gat,s3083gat,s609gat);
  nor x1043(s3147gat,s2930gat,s3083gat);
  nor x1044(s3150gat,s3034gat,s3087gat);
  nor x1045(s3151gat,s3087gat,s657gat);
  nor x1046(s3152gat,s2934gat,s3087gat);
  nor x1047(s3155gat,s3037gat,s3091gat);
  nor x1048(s3156gat,s3091gat,s705gat);
  nor x1049(s3157gat,s2938gat,s3091gat);
  nor x1050(s3160gat,s3040gat,s3095gat);
  nor x1051(s3161gat,s3095gat,s753gat);
  nor x1052(s3162gat,s2942gat,s3095gat);
  nor x1053(s3165gat,s3043gat,s3099gat);
  nor x1054(s3166gat,s3099gat,s801gat);
  nor x1055(s3167gat,s2946gat,s3099gat);
  nor x1056(s3170gat,s3046gat,s3103gat);
  nor x1057(s3171gat,s3103gat,s849gat);
  nor x1058(s3172gat,s2950gat,s3103gat);
  nor x1059(s3175gat,s3049gat,s3107gat);
  nor x1060(s3176gat,s3107gat,s897gat);
  nor x1061(s3177gat,s2954gat,s3107gat);
  nor x1062(s3180gat,s3052gat,s3111gat);
  nor x1063(s3181gat,s3111gat,s945gat);
  nor x1064(s3182gat,s2958gat,s3111gat);
  nor x1065(s3185gat,s3055gat,s3115gat);
  nor x1066(s3186gat,s3115gat,s993gat);
  nor x1067(s3187gat,s2962gat,s3115gat);
  nor x1068(s3190gat,s3119gat,s3120gat);
  nor x1069(s3193gat,s3124gat,s3121gat);
  nor x1070(s3197gat,s3067gat,s3127gat);
  nor x1071(s3198gat,s3127gat,s3064gat);
  nor x1072(s3199gat,s3131gat,s3132gat);
  nor x1073(s3202gat,s3133gat,s1188gat);
  nor x1074(s3206gat,s3076gat,s3136gat);
  nor x1075(s3207gat,s3136gat,s1236gat);
  nor x1076(s3208gat,s2983gat,s3136gat);
  nor x1077(s3211gat,s3140gat,s3141gat);
  nor x1078(s3212gat,s3145gat,s3146gat);
  nor x1079(s3215gat,s3150gat,s3151gat);
  nor x1080(s3218gat,s3155gat,s3156gat);
  nor x1081(s3221gat,s3160gat,s3161gat);
  nor x1082(s3224gat,s3165gat,s3166gat);
  nor x1083(s3227gat,s3170gat,s3171gat);
  nor x1084(s3230gat,s3175gat,s3176gat);
  nor x1085(s3233gat,s3180gat,s3181gat);
  nor x1086(s3236gat,s3185gat,s3186gat);
  nor x1087(s3239gat,s3190gat,s3187gat);
  nor x1088(s3243gat,s3124gat,s3193gat);
  nor x1089(s3244gat,s3193gat,s3121gat);
  nor x1090(s3245gat,s3197gat,s3198gat);
  nor x1091(s3248gat,s3199gat,s1140gat);
  nor x1092(s3252gat,s3133gat,s3202gat);
  nor x1093(s3253gat,s3202gat,s1188gat);
  nor x1094(s3254gat,s3022gat,s3202gat);
  nor x1095(s3257gat,s3206gat,s3207gat);
  nor x1096(s3260gat,s1284gat,s3208gat);
  nor x1097(s3264gat,s3212gat,s3142gat);
  nor x1098(s3268gat,s3215gat,s3147gat);
  nor x1099(s3272gat,s3218gat,s3152gat);
  nor x1100(s3276gat,s3221gat,s3157gat);
  nor x1101(s3280gat,s3224gat,s3162gat);
  nor x1102(s3284gat,s3227gat,s3167gat);
  nor x1103(s3288gat,s3230gat,s3172gat);
  nor x1104(s3292gat,s3233gat,s3177gat);
  nor x1105(s3296gat,s3236gat,s3182gat);
  nor x1106(s3300gat,s3190gat,s3239gat);
  nor x1107(s3301gat,s3239gat,s3187gat);
  nor x1108(s3302gat,s3243gat,s3244gat);
  nor x1109(s3305gat,s3245gat,s1092gat);
  nor x1110(s3309gat,s3199gat,s3248gat);
  nor x1111(s3310gat,s3248gat,s1140gat);
  nor x1112(s3311gat,s3070gat,s3248gat);
  nor x1113(s3314gat,s3252gat,s3253gat);
  nor x1114(s3317gat,s3257gat,s3254gat);
  nor x1115(s3321gat,s1284gat,s3260gat);
  nor x1116(s3322gat,s3260gat,s3208gat);
  nor x1117(s3323gat,s3212gat,s3264gat);
  nor x1118(s3324gat,s3264gat,s3142gat);
  nor x1119(s3325gat,s3215gat,s3268gat);
  nor x1120(s3326gat,s3268gat,s3147gat);
  nor x1121(s3327gat,s3218gat,s3272gat);
  nor x1122(s3328gat,s3272gat,s3152gat);
  nor x1123(s3329gat,s3221gat,s3276gat);
  nor x1124(s3330gat,s3276gat,s3157gat);
  nor x1125(s3331gat,s3224gat,s3280gat);
  nor x1126(s3332gat,s3280gat,s3162gat);
  nor x1127(s3333gat,s3227gat,s3284gat);
  nor x1128(s3334gat,s3284gat,s3167gat);
  nor x1129(s3335gat,s3230gat,s3288gat);
  nor x1130(s3336gat,s3288gat,s3172gat);
  nor x1131(s3337gat,s3233gat,s3292gat);
  nor x1132(s3338gat,s3292gat,s3177gat);
  nor x1133(s3339gat,s3236gat,s3296gat);
  nor x1134(s3340gat,s3296gat,s3182gat);
  nor x1135(s3341gat,s3300gat,s3301gat);
  nor x1136(s3344gat,s3302gat,s1044gat);
  nor x1137(s3348gat,s3245gat,s3305gat);
  nor x1138(s3349gat,s3305gat,s1092gat);
  nor x1139(s3350gat,s3127gat,s3305gat);
  nor x1140(s3353gat,s3309gat,s3310gat);
  nor x1141(s3356gat,s3314gat,s3311gat);
  nor x1142(s3360gat,s3257gat,s3317gat);
  nor x1143(s3361gat,s3317gat,s3254gat);
  nor x1144(s3362gat,s3321gat,s3322gat);
  nor x1145(s3365gat,s3323gat,s3324gat);
  nor x1146(s3368gat,s3325gat,s3326gat);
  nor x1147(s3371gat,s3327gat,s3328gat);
  nor x1148(s3374gat,s3329gat,s3330gat);
  nor x1149(s3377gat,s3331gat,s3332gat);
  nor x1150(s3380gat,s3333gat,s3334gat);
  nor x1151(s3383gat,s3335gat,s3336gat);
  nor x1152(s3386gat,s3337gat,s3338gat);
  nor x1153(s3389gat,s3339gat,s3340gat);
  nor x1154(s3392gat,s3341gat,s996gat);
  nor x1155(s3396gat,s3302gat,s3344gat);
  nor x1156(s3397gat,s3344gat,s1044gat);
  nor x1157(s3398gat,s3193gat,s3344gat);
  nor x1158(s3401gat,s3348gat,s3349gat);
  nor x1159(s3404gat,s3353gat,s3350gat);
  nor x1160(s3408gat,s3314gat,s3356gat);
  nor x1161(s3409gat,s3356gat,s3311gat);
  nor x1162(s3410gat,s3360gat,s3361gat);
  nor x1163(s3413gat,s3362gat,s1239gat);
  nor x1164(s3417gat,s3365gat,s564gat);
  nor x1165(s3421gat,s3368gat,s612gat);
  nor x1166(s3425gat,s3371gat,s660gat);
  nor x1167(s3429gat,s3374gat,s708gat);
  nor x1168(s3433gat,s3377gat,s756gat);
  nor x1169(s3437gat,s3380gat,s804gat);
  nor x1170(s3441gat,s3383gat,s852gat);
  nor x1171(s3445gat,s3386gat,s900gat);
  nor x1172(s3449gat,s3389gat,s948gat);
  nor x1173(s3453gat,s3341gat,s3392gat);
  nor x1174(s3454gat,s3392gat,s996gat);
  nor x1175(s3455gat,s3239gat,s3392gat);
  nor x1176(s3458gat,s3396gat,s3397gat);
  nor x1177(s3461gat,s3401gat,s3398gat);
  nor x1178(s3465gat,s3353gat,s3404gat);
  nor x1179(s3466gat,s3404gat,s3350gat);
  nor x1180(s3467gat,s3408gat,s3409gat);
  nor x1181(s3470gat,s3410gat,s1191gat);
  nor x1182(s3474gat,s3362gat,s3413gat);
  nor x1183(s3475gat,s3413gat,s1239gat);
  nor x1184(s3476gat,s3260gat,s3413gat);
  nor x1185(s3479gat,s3365gat,s3417gat);
  nor x1186(s3480gat,s3417gat,s564gat);
  nor x1187(s3481gat,s3264gat,s3417gat);
  nor x1188(s3484gat,s3368gat,s3421gat);
  nor x1189(s3485gat,s3421gat,s612gat);
  nor x1190(s3486gat,s3268gat,s3421gat);
  nor x1191(s3489gat,s3371gat,s3425gat);
  nor x1192(s3490gat,s3425gat,s660gat);
  nor x1193(s3491gat,s3272gat,s3425gat);
  nor x1194(s3494gat,s3374gat,s3429gat);
  nor x1195(s3495gat,s3429gat,s708gat);
  nor x1196(s3496gat,s3276gat,s3429gat);
  nor x1197(s3499gat,s3377gat,s3433gat);
  nor x1198(s3500gat,s3433gat,s756gat);
  nor x1199(s3501gat,s3280gat,s3433gat);
  nor x1200(s3504gat,s3380gat,s3437gat);
  nor x1201(s3505gat,s3437gat,s804gat);
  nor x1202(s3506gat,s3284gat,s3437gat);
  nor x1203(s3509gat,s3383gat,s3441gat);
  nor x1204(s3510gat,s3441gat,s852gat);
  nor x1205(s3511gat,s3288gat,s3441gat);
  nor x1206(s3514gat,s3386gat,s3445gat);
  nor x1207(s3515gat,s3445gat,s900gat);
  nor x1208(s3516gat,s3292gat,s3445gat);
  nor x1209(s3519gat,s3389gat,s3449gat);
  nor x1210(s3520gat,s3449gat,s948gat);
  nor x1211(s3521gat,s3296gat,s3449gat);
  nor x1212(s3524gat,s3453gat,s3454gat);
  nor x1213(s3527gat,s3458gat,s3455gat);
  nor x1214(s3531gat,s3401gat,s3461gat);
  nor x1215(s3532gat,s3461gat,s3398gat);
  nor x1216(s3533gat,s3465gat,s3466gat);
  nor x1217(s3536gat,s3467gat,s1143gat);
  nor x1218(s3540gat,s3410gat,s3470gat);
  nor x1219(s3541gat,s3470gat,s1191gat);
  nor x1220(s3542gat,s3317gat,s3470gat);
  nor x1221(s3545gat,s3474gat,s3475gat);
  nor x1222(s3548gat,s1287gat,s3476gat);
  nor x1223(s3552gat,s3479gat,s3480gat);
  nor x1224(s3553gat,s3484gat,s3485gat);
  nor x1225(s3556gat,s3489gat,s3490gat);
  nor x1226(s3559gat,s3494gat,s3495gat);
  nor x1227(s3562gat,s3499gat,s3500gat);
  nor x1228(s3565gat,s3504gat,s3505gat);
  nor x1229(s3568gat,s3509gat,s3510gat);
  nor x1230(s3571gat,s3514gat,s3515gat);
  nor x1231(s3574gat,s3519gat,s3520gat);
  nor x1232(s3577gat,s3524gat,s3521gat);
  nor x1233(s3581gat,s3458gat,s3527gat);
  nor x1234(s3582gat,s3527gat,s3455gat);
  nor x1235(s3583gat,s3531gat,s3532gat);
  nor x1236(s3586gat,s3533gat,s1095gat);
  nor x1237(s3590gat,s3467gat,s3536gat);
  nor x1238(s3591gat,s3536gat,s1143gat);
  nor x1239(s3592gat,s3356gat,s3536gat);
  nor x1240(s3595gat,s3540gat,s3541gat);
  nor x1241(s3598gat,s3545gat,s3542gat);
  nor x1242(s3602gat,s1287gat,s3548gat);
  nor x1243(s3603gat,s3548gat,s3476gat);
  nor x1244(s3604gat,s3553gat,s3481gat);
  nor x1245(s3608gat,s3556gat,s3486gat);
  nor x1246(s3612gat,s3559gat,s3491gat);
  nor x1247(s3616gat,s3562gat,s3496gat);
  nor x1248(s3620gat,s3565gat,s3501gat);
  nor x1249(s3624gat,s3568gat,s3506gat);
  nor x1250(s3628gat,s3571gat,s3511gat);
  nor x1251(s3632gat,s3574gat,s3516gat);
  nor x1252(s3636gat,s3524gat,s3577gat);
  nor x1253(s3637gat,s3577gat,s3521gat);
  nor x1254(s3638gat,s3581gat,s3582gat);
  nor x1255(s3641gat,s3583gat,s1047gat);
  nor x1256(s3645gat,s3533gat,s3586gat);
  nor x1257(s3646gat,s3586gat,s1095gat);
  nor x1258(s3647gat,s3404gat,s3586gat);
  nor x1259(s3650gat,s3590gat,s3591gat);
  nor x1260(s3653gat,s3595gat,s3592gat);
  nor x1261(s3657gat,s3545gat,s3598gat);
  nor x1262(s3658gat,s3598gat,s3542gat);
  nor x1263(s3659gat,s3602gat,s3603gat);
  nor x1264(s3662gat,s3553gat,s3604gat);
  nor x1265(s3663gat,s3604gat,s3481gat);
  nor x1266(s3664gat,s3556gat,s3608gat);
  nor x1267(s3665gat,s3608gat,s3486gat);
  nor x1268(s3666gat,s3559gat,s3612gat);
  nor x1269(s3667gat,s3612gat,s3491gat);
  nor x1270(s3668gat,s3562gat,s3616gat);
  nor x1271(s3669gat,s3616gat,s3496gat);
  nor x1272(s3670gat,s3565gat,s3620gat);
  nor x1273(s3671gat,s3620gat,s3501gat);
  nor x1274(s3672gat,s3568gat,s3624gat);
  nor x1275(s3673gat,s3624gat,s3506gat);
  nor x1276(s3674gat,s3571gat,s3628gat);
  nor x1277(s3675gat,s3628gat,s3511gat);
  nor x1278(s3676gat,s3574gat,s3632gat);
  nor x1279(s3677gat,s3632gat,s3516gat);
  nor x1280(s3678gat,s3636gat,s3637gat);
  nor x1281(s3681gat,s3638gat,s999gat);
  nor x1282(s3685gat,s3583gat,s3641gat);
  nor x1283(s3686gat,s3641gat,s1047gat);
  nor x1284(s3687gat,s3461gat,s3641gat);
  nor x1285(s3690gat,s3645gat,s3646gat);
  nor x1286(s3693gat,s3650gat,s3647gat);
  nor x1287(s3697gat,s3595gat,s3653gat);
  nor x1288(s3698gat,s3653gat,s3592gat);
  nor x1289(s3699gat,s3657gat,s3658gat);
  nor x1290(s3702gat,s3659gat,s1242gat);
  nor x1291(s3706gat,s3662gat,s3663gat);
  nor x1292(s3709gat,s3664gat,s3665gat);
  nor x1293(s3712gat,s3666gat,s3667gat);
  nor x1294(s3715gat,s3668gat,s3669gat);
  nor x1295(s3718gat,s3670gat,s3671gat);
  nor x1296(s3721gat,s3672gat,s3673gat);
  nor x1297(s3724gat,s3674gat,s3675gat);
  nor x1298(s3727gat,s3676gat,s3677gat);
  nor x1299(s3730gat,s3678gat,s951gat);
  nor x1300(s3734gat,s3638gat,s3681gat);
  nor x1301(s3735gat,s3681gat,s999gat);
  nor x1302(s3736gat,s3527gat,s3681gat);
  nor x1303(s3739gat,s3685gat,s3686gat);
  nor x1304(s3742gat,s3690gat,s3687gat);
  nor x1305(s3746gat,s3650gat,s3693gat);
  nor x1306(s3747gat,s3693gat,s3647gat);
  nor x1307(s3748gat,s3697gat,s3698gat);
  nor x1308(s3751gat,s3699gat,s1194gat);
  nor x1309(s3755gat,s3659gat,s3702gat);
  nor x1310(s3756gat,s3702gat,s1242gat);
  nor x1311(s3757gat,s3548gat,s3702gat);
  nor x1312(s3760gat,s3706gat,s567gat);
  nor x1313(s3764gat,s3709gat,s615gat);
  nor x1314(s3768gat,s3712gat,s663gat);
  nor x1315(s3772gat,s3715gat,s711gat);
  nor x1316(s3776gat,s3718gat,s759gat);
  nor x1317(s3780gat,s3721gat,s807gat);
  nor x1318(s3784gat,s3724gat,s855gat);
  nor x1319(s3788gat,s3727gat,s903gat);
  nor x1320(s3792gat,s3678gat,s3730gat);
  nor x1321(s3793gat,s3730gat,s951gat);
  nor x1322(s3794gat,s3577gat,s3730gat);
  nor x1323(s3797gat,s3734gat,s3735gat);
  nor x1324(s3800gat,s3739gat,s3736gat);
  nor x1325(s3804gat,s3690gat,s3742gat);
  nor x1326(s3805gat,s3742gat,s3687gat);
  nor x1327(s3806gat,s3746gat,s3747gat);
  nor x1328(s3809gat,s3748gat,s1146gat);
  nor x1329(s3813gat,s3699gat,s3751gat);
  nor x1330(s3814gat,s3751gat,s1194gat);
  nor x1331(s3815gat,s3598gat,s3751gat);
  nor x1332(s3818gat,s3755gat,s3756gat);
  nor x1333(s3821gat,s1290gat,s3757gat);
  nor x1334(s3825gat,s3706gat,s3760gat);
  nor x1335(s3826gat,s3760gat,s567gat);
  nor x1336(s3827gat,s3604gat,s3760gat);
  nor x1337(s3830gat,s3709gat,s3764gat);
  nor x1338(s3831gat,s3764gat,s615gat);
  nor x1339(s3832gat,s3608gat,s3764gat);
  nor x1340(s3835gat,s3712gat,s3768gat);
  nor x1341(s3836gat,s3768gat,s663gat);
  nor x1342(s3837gat,s3612gat,s3768gat);
  nor x1343(s3840gat,s3715gat,s3772gat);
  nor x1344(s3841gat,s3772gat,s711gat);
  nor x1345(s3842gat,s3616gat,s3772gat);
  nor x1346(s3845gat,s3718gat,s3776gat);
  nor x1347(s3846gat,s3776gat,s759gat);
  nor x1348(s3847gat,s3620gat,s3776gat);
  nor x1349(s3850gat,s3721gat,s3780gat);
  nor x1350(s3851gat,s3780gat,s807gat);
  nor x1351(s3852gat,s3624gat,s3780gat);
  nor x1352(s3855gat,s3724gat,s3784gat);
  nor x1353(s3856gat,s3784gat,s855gat);
  nor x1354(s3857gat,s3628gat,s3784gat);
  nor x1355(s3860gat,s3727gat,s3788gat);
  nor x1356(s3861gat,s3788gat,s903gat);
  nor x1357(s3862gat,s3632gat,s3788gat);
  nor x1358(s3865gat,s3792gat,s3793gat);
  nor x1359(s3868gat,s3797gat,s3794gat);
  nor x1360(s3872gat,s3739gat,s3800gat);
  nor x1361(s3873gat,s3800gat,s3736gat);
  nor x1362(s3874gat,s3804gat,s3805gat);
  nor x1363(s3877gat,s3806gat,s1098gat);
  nor x1364(s3881gat,s3748gat,s3809gat);
  nor x1365(s3882gat,s3809gat,s1146gat);
  nor x1366(s3883gat,s3653gat,s3809gat);
  nor x1367(s3886gat,s3813gat,s3814gat);
  nor x1368(s3889gat,s3818gat,s3815gat);
  nor x1369(s3893gat,s1290gat,s3821gat);
  nor x1370(s3894gat,s3821gat,s3757gat);
  nor x1371(s3895gat,s3825gat,s3826gat);
  nor x1372(s3896gat,s3830gat,s3831gat);
  nor x1373(s3899gat,s3835gat,s3836gat);
  nor x1374(s3902gat,s3840gat,s3841gat);
  nor x1375(s3905gat,s3845gat,s3846gat);
  nor x1376(s3908gat,s3850gat,s3851gat);
  nor x1377(s3911gat,s3855gat,s3856gat);
  nor x1378(s3914gat,s3860gat,s3861gat);
  nor x1379(s3917gat,s3865gat,s3862gat);
  nor x1380(s3921gat,s3797gat,s3868gat);
  nor x1381(s3922gat,s3868gat,s3794gat);
  nor x1382(s3923gat,s3872gat,s3873gat);
  nor x1383(s3926gat,s3874gat,s1050gat);
  nor x1384(s3930gat,s3806gat,s3877gat);
  nor x1385(s3931gat,s3877gat,s1098gat);
  nor x1386(s3932gat,s3693gat,s3877gat);
  nor x1387(s3935gat,s3881gat,s3882gat);
  nor x1388(s3938gat,s3886gat,s3883gat);
  nor x1389(s3942gat,s3818gat,s3889gat);
  nor x1390(s3943gat,s3889gat,s3815gat);
  nor x1391(s3944gat,s3893gat,s3894gat);
  nor x1392(s3947gat,s3896gat,s3827gat);
  nor x1393(s3951gat,s3899gat,s3832gat);
  nor x1394(s3955gat,s3902gat,s3837gat);
  nor x1395(s3959gat,s3905gat,s3842gat);
  nor x1396(s3963gat,s3908gat,s3847gat);
  nor x1397(s3967gat,s3911gat,s3852gat);
  nor x1398(s3971gat,s3914gat,s3857gat);
  nor x1399(s3975gat,s3865gat,s3917gat);
  nor x1400(s3976gat,s3917gat,s3862gat);
  nor x1401(s3977gat,s3921gat,s3922gat);
  nor x1402(s3980gat,s3923gat,s1002gat);
  nor x1403(s3984gat,s3874gat,s3926gat);
  nor x1404(s3985gat,s3926gat,s1050gat);
  nor x1405(s3986gat,s3742gat,s3926gat);
  nor x1406(s3989gat,s3930gat,s3931gat);
  nor x1407(s3992gat,s3935gat,s3932gat);
  nor x1408(s3996gat,s3886gat,s3938gat);
  nor x1409(s3997gat,s3938gat,s3883gat);
  nor x1410(s3998gat,s3942gat,s3943gat);
  nor x1411(s4001gat,s3944gat,s1245gat);
  nor x1412(s4005gat,s3896gat,s3947gat);
  nor x1413(s4006gat,s3947gat,s3827gat);
  nor x1414(s4007gat,s3899gat,s3951gat);
  nor x1415(s4008gat,s3951gat,s3832gat);
  nor x1416(s4009gat,s3902gat,s3955gat);
  nor x1417(s4010gat,s3955gat,s3837gat);
  nor x1418(s4011gat,s3905gat,s3959gat);
  nor x1419(s4012gat,s3959gat,s3842gat);
  nor x1420(s4013gat,s3908gat,s3963gat);
  nor x1421(s4014gat,s3963gat,s3847gat);
  nor x1422(s4015gat,s3911gat,s3967gat);
  nor x1423(s4016gat,s3967gat,s3852gat);
  nor x1424(s4017gat,s3914gat,s3971gat);
  nor x1425(s4018gat,s3971gat,s3857gat);
  nor x1426(s4019gat,s3975gat,s3976gat);
  nor x1427(s4022gat,s3977gat,s954gat);
  nor x1428(s4026gat,s3923gat,s3980gat);
  nor x1429(s4027gat,s3980gat,s1002gat);
  nor x1430(s4028gat,s3800gat,s3980gat);
  nor x1431(s4031gat,s3984gat,s3985gat);
  nor x1432(s4034gat,s3989gat,s3986gat);
  nor x1433(s4038gat,s3935gat,s3992gat);
  nor x1434(s4039gat,s3992gat,s3932gat);
  nor x1435(s4040gat,s3996gat,s3997gat);
  nor x1436(s4043gat,s3998gat,s1197gat);
  nor x1437(s4047gat,s3944gat,s4001gat);
  nor x1438(s4048gat,s4001gat,s1245gat);
  nor x1439(s4049gat,s3821gat,s4001gat);
  nor x1440(s4052gat,s4005gat,s4006gat);
  nor x1441(s4055gat,s4007gat,s4008gat);
  nor x1442(s4058gat,s4009gat,s4010gat);
  nor x1443(s4061gat,s4011gat,s4012gat);
  nor x1444(s4064gat,s4013gat,s4014gat);
  nor x1445(s4067gat,s4015gat,s4016gat);
  nor x1446(s4070gat,s4017gat,s4018gat);
  nor x1447(s4073gat,s4019gat,s906gat);
  nor x1448(s4077gat,s3977gat,s4022gat);
  nor x1449(s4078gat,s4022gat,s954gat);
  nor x1450(s4079gat,s3868gat,s4022gat);
  nor x1451(s4082gat,s4026gat,s4027gat);
  nor x1452(s4085gat,s4031gat,s4028gat);
  nor x1453(s4089gat,s3989gat,s4034gat);
  nor x1454(s4090gat,s4034gat,s3986gat);
  nor x1455(s4091gat,s4038gat,s4039gat);
  nor x1456(s4094gat,s4040gat,s1149gat);
  nor x1457(s4098gat,s3998gat,s4043gat);
  nor x1458(s4099gat,s4043gat,s1197gat);
  nor x1459(s4100gat,s3889gat,s4043gat);
  nor x1460(s4103gat,s4047gat,s4048gat);
  nor x1461(s4106gat,s1293gat,s4049gat);
  nor x1462(s4110gat,s4052gat,s570gat);
  nor x1463(s4114gat,s4055gat,s618gat);
  nor x1464(s4118gat,s4058gat,s666gat);
  nor x1465(s4122gat,s4061gat,s714gat);
  nor x1466(s4126gat,s4064gat,s762gat);
  nor x1467(s4130gat,s4067gat,s810gat);
  nor x1468(s4134gat,s4070gat,s858gat);
  nor x1469(s4138gat,s4019gat,s4073gat);
  nor x1470(s4139gat,s4073gat,s906gat);
  nor x1471(s4140gat,s3917gat,s4073gat);
  nor x1472(s4143gat,s4077gat,s4078gat);
  nor x1473(s4146gat,s4082gat,s4079gat);
  nor x1474(s4150gat,s4031gat,s4085gat);
  nor x1475(s4151gat,s4085gat,s4028gat);
  nor x1476(s4152gat,s4089gat,s4090gat);
  nor x1477(s4155gat,s4091gat,s1101gat);
  nor x1478(s4159gat,s4040gat,s4094gat);
  nor x1479(s4160gat,s4094gat,s1149gat);
  nor x1480(s4161gat,s3938gat,s4094gat);
  nor x1481(s4164gat,s4098gat,s4099gat);
  nor x1482(s4167gat,s4103gat,s4100gat);
  nor x1483(s4171gat,s1293gat,s4106gat);
  nor x1484(s4172gat,s4106gat,s4049gat);
  nor x1485(s4173gat,s4052gat,s4110gat);
  nor x1486(s4174gat,s4110gat,s570gat);
  nor x1487(s4175gat,s3947gat,s4110gat);
  nor x1488(s4178gat,s4055gat,s4114gat);
  nor x1489(s4179gat,s4114gat,s618gat);
  nor x1490(s4180gat,s3951gat,s4114gat);
  nor x1491(s4183gat,s4058gat,s4118gat);
  nor x1492(s4184gat,s4118gat,s666gat);
  nor x1493(s4185gat,s3955gat,s4118gat);
  nor x1494(s4188gat,s4061gat,s4122gat);
  nor x1495(s4189gat,s4122gat,s714gat);
  nor x1496(s4190gat,s3959gat,s4122gat);
  nor x1497(s4193gat,s4064gat,s4126gat);
  nor x1498(s4194gat,s4126gat,s762gat);
  nor x1499(s4195gat,s3963gat,s4126gat);
  nor x1500(s4198gat,s4067gat,s4130gat);
  nor x1501(s4199gat,s4130gat,s810gat);
  nor x1502(s4200gat,s3967gat,s4130gat);
  nor x1503(s4203gat,s4070gat,s4134gat);
  nor x1504(s4204gat,s4134gat,s858gat);
  nor x1505(s4205gat,s3971gat,s4134gat);
  nor x1506(s4208gat,s4138gat,s4139gat);
  nor x1507(s4211gat,s4143gat,s4140gat);
  nor x1508(s4215gat,s4082gat,s4146gat);
  nor x1509(s4216gat,s4146gat,s4079gat);
  nor x1510(s4217gat,s4150gat,s4151gat);
  nor x1511(s4220gat,s4152gat,s1053gat);
  nor x1512(s4224gat,s4091gat,s4155gat);
  nor x1513(s4225gat,s4155gat,s1101gat);
  nor x1514(s4226gat,s3992gat,s4155gat);
  nor x1515(s4229gat,s4159gat,s4160gat);
  nor x1516(s4232gat,s4164gat,s4161gat);
  nor x1517(s4236gat,s4103gat,s4167gat);
  nor x1518(s4237gat,s4167gat,s4100gat);
  nor x1519(s4238gat,s4171gat,s4172gat);
  nor x1520(s4241gat,s4173gat,s4174gat);
  nor x1521(s4242gat,s4178gat,s4179gat);
  nor x1522(s4245gat,s4183gat,s4184gat);
  nor x1523(s4248gat,s4188gat,s4189gat);
  nor x1524(s4251gat,s4193gat,s4194gat);
  nor x1525(s4254gat,s4198gat,s4199gat);
  nor x1526(s4257gat,s4203gat,s4204gat);
  nor x1527(s4260gat,s4208gat,s4205gat);
  nor x1528(s4264gat,s4143gat,s4211gat);
  nor x1529(s4265gat,s4211gat,s4140gat);
  nor x1530(s4266gat,s4215gat,s4216gat);
  nor x1531(s4269gat,s4217gat,s1005gat);
  nor x1532(s4273gat,s4152gat,s4220gat);
  nor x1533(s4274gat,s4220gat,s1053gat);
  nor x1534(s4275gat,s4034gat,s4220gat);
  nor x1535(s4278gat,s4224gat,s4225gat);
  nor x1536(s4281gat,s4229gat,s4226gat);
  nor x1537(s4285gat,s4164gat,s4232gat);
  nor x1538(s4286gat,s4232gat,s4161gat);
  nor x1539(s4287gat,s4236gat,s4237gat);
  nor x1540(s4290gat,s4238gat,s1248gat);
  nor x1541(s4294gat,s4242gat,s4175gat);
  nor x1542(s4298gat,s4245gat,s4180gat);
  nor x1543(s4302gat,s4248gat,s4185gat);
  nor x1544(s4306gat,s4251gat,s4190gat);
  nor x1545(s4310gat,s4254gat,s4195gat);
  nor x1546(s4314gat,s4257gat,s4200gat);
  nor x1547(s4318gat,s4208gat,s4260gat);
  nor x1548(s4319gat,s4260gat,s4205gat);
  nor x1549(s4320gat,s4264gat,s4265gat);
  nor x1550(s4323gat,s4266gat,s957gat);
  nor x1551(s4327gat,s4217gat,s4269gat);
  nor x1552(s4328gat,s4269gat,s1005gat);
  nor x1553(s4329gat,s4085gat,s4269gat);
  nor x1554(s4332gat,s4273gat,s4274gat);
  nor x1555(s4335gat,s4278gat,s4275gat);
  nor x1556(s4339gat,s4229gat,s4281gat);
  nor x1557(s4340gat,s4281gat,s4226gat);
  nor x1558(s4341gat,s4285gat,s4286gat);
  nor x1559(s4344gat,s4287gat,s1200gat);
  nor x1560(s4348gat,s4238gat,s4290gat);
  nor x1561(s4349gat,s4290gat,s1248gat);
  nor x1562(s4350gat,s4106gat,s4290gat);
  nor x1563(s4353gat,s4242gat,s4294gat);
  nor x1564(s4354gat,s4294gat,s4175gat);
  nor x1565(s4355gat,s4245gat,s4298gat);
  nor x1566(s4356gat,s4298gat,s4180gat);
  nor x1567(s4357gat,s4248gat,s4302gat);
  nor x1568(s4358gat,s4302gat,s4185gat);
  nor x1569(s4359gat,s4251gat,s4306gat);
  nor x1570(s4360gat,s4306gat,s4190gat);
  nor x1571(s4361gat,s4254gat,s4310gat);
  nor x1572(s4362gat,s4310gat,s4195gat);
  nor x1573(s4363gat,s4257gat,s4314gat);
  nor x1574(s4364gat,s4314gat,s4200gat);
  nor x1575(s4365gat,s4318gat,s4319gat);
  nor x1576(s4368gat,s4320gat,s909gat);
  nor x1577(s4372gat,s4266gat,s4323gat);
  nor x1578(s4373gat,s4323gat,s957gat);
  nor x1579(s4374gat,s4146gat,s4323gat);
  nor x1580(s4377gat,s4327gat,s4328gat);
  nor x1581(s4380gat,s4332gat,s4329gat);
  nor x1582(s4384gat,s4278gat,s4335gat);
  nor x1583(s4385gat,s4335gat,s4275gat);
  nor x1584(s4386gat,s4339gat,s4340gat);
  nor x1585(s4389gat,s4341gat,s1152gat);
  nor x1586(s4393gat,s4287gat,s4344gat);
  nor x1587(s4394gat,s4344gat,s1200gat);
  nor x1588(s4395gat,s4167gat,s4344gat);
  nor x1589(s4398gat,s4348gat,s4349gat);
  nor x1590(s4401gat,s1296gat,s4350gat);
  nor x1591(s4405gat,s4353gat,s4354gat);
  nor x1592(s4408gat,s4355gat,s4356gat);
  nor x1593(s4411gat,s4357gat,s4358gat);
  nor x1594(s4414gat,s4359gat,s4360gat);
  nor x1595(s4417gat,s4361gat,s4362gat);
  nor x1596(s4420gat,s4363gat,s4364gat);
  nor x1597(s4423gat,s4365gat,s861gat);
  nor x1598(s4427gat,s4320gat,s4368gat);
  nor x1599(s4428gat,s4368gat,s909gat);
  nor x1600(s4429gat,s4211gat,s4368gat);
  nor x1601(s4432gat,s4372gat,s4373gat);
  nor x1602(s4435gat,s4377gat,s4374gat);
  nor x1603(s4439gat,s4332gat,s4380gat);
  nor x1604(s4440gat,s4380gat,s4329gat);
  nor x1605(s4441gat,s4384gat,s4385gat);
  nor x1606(s4444gat,s4386gat,s1104gat);
  nor x1607(s4448gat,s4341gat,s4389gat);
  nor x1608(s4449gat,s4389gat,s1152gat);
  nor x1609(s4450gat,s4232gat,s4389gat);
  nor x1610(s4453gat,s4393gat,s4394gat);
  nor x1611(s4456gat,s4398gat,s4395gat);
  nor x1612(s4460gat,s1296gat,s4401gat);
  nor x1613(s4461gat,s4401gat,s4350gat);
  nor x1614(s4462gat,s4405gat,s573gat);
  nor x1615(s4466gat,s4408gat,s621gat);
  nor x1616(s4470gat,s4411gat,s669gat);
  nor x1617(s4474gat,s4414gat,s717gat);
  nor x1618(s4478gat,s4417gat,s765gat);
  nor x1619(s4482gat,s4420gat,s813gat);
  nor x1620(s4486gat,s4365gat,s4423gat);
  nor x1621(s4487gat,s4423gat,s861gat);
  nor x1622(s4488gat,s4260gat,s4423gat);
  nor x1623(s4491gat,s4427gat,s4428gat);
  nor x1624(s4494gat,s4432gat,s4429gat);
  nor x1625(s4498gat,s4377gat,s4435gat);
  nor x1626(s4499gat,s4435gat,s4374gat);
  nor x1627(s4500gat,s4439gat,s4440gat);
  nor x1628(s4503gat,s4441gat,s1056gat);
  nor x1629(s4507gat,s4386gat,s4444gat);
  nor x1630(s4508gat,s4444gat,s1104gat);
  nor x1631(s4509gat,s4281gat,s4444gat);
  nor x1632(s4512gat,s4448gat,s4449gat);
  nor x1633(s4515gat,s4453gat,s4450gat);
  nor x1634(s4519gat,s4398gat,s4456gat);
  nor x1635(s4520gat,s4456gat,s4395gat);
  nor x1636(s4521gat,s4460gat,s4461gat);
  nor x1637(s4524gat,s4405gat,s4462gat);
  nor x1638(s4525gat,s4462gat,s573gat);
  nor x1639(s4526gat,s4294gat,s4462gat);
  nor x1640(s4529gat,s4408gat,s4466gat);
  nor x1641(s4530gat,s4466gat,s621gat);
  nor x1642(s4531gat,s4298gat,s4466gat);
  nor x1643(s4534gat,s4411gat,s4470gat);
  nor x1644(s4535gat,s4470gat,s669gat);
  nor x1645(s4536gat,s4302gat,s4470gat);
  nor x1646(s4539gat,s4414gat,s4474gat);
  nor x1647(s4540gat,s4474gat,s717gat);
  nor x1648(s4541gat,s4306gat,s4474gat);
  nor x1649(s4544gat,s4417gat,s4478gat);
  nor x1650(s4545gat,s4478gat,s765gat);
  nor x1651(s4546gat,s4310gat,s4478gat);
  nor x1652(s4549gat,s4420gat,s4482gat);
  nor x1653(s4550gat,s4482gat,s813gat);
  nor x1654(s4551gat,s4314gat,s4482gat);
  nor x1655(s4554gat,s4486gat,s4487gat);
  nor x1656(s4557gat,s4491gat,s4488gat);
  nor x1657(s4561gat,s4432gat,s4494gat);
  nor x1658(s4562gat,s4494gat,s4429gat);
  nor x1659(s4563gat,s4498gat,s4499gat);
  nor x1660(s4566gat,s4500gat,s1008gat);
  nor x1661(s4570gat,s4441gat,s4503gat);
  nor x1662(s4571gat,s4503gat,s1056gat);
  nor x1663(s4572gat,s4335gat,s4503gat);
  nor x1664(s4575gat,s4507gat,s4508gat);
  nor x1665(s4578gat,s4512gat,s4509gat);
  nor x1666(s4582gat,s4453gat,s4515gat);
  nor x1667(s4583gat,s4515gat,s4450gat);
  nor x1668(s4584gat,s4519gat,s4520gat);
  nor x1669(s4587gat,s4521gat,s1251gat);
  nor x1670(s4591gat,s4524gat,s4525gat);
  nor x1671(s4592gat,s4529gat,s4530gat);
  nor x1672(s4595gat,s4534gat,s4535gat);
  nor x1673(s4598gat,s4539gat,s4540gat);
  nor x1674(s4601gat,s4544gat,s4545gat);
  nor x1675(s4604gat,s4549gat,s4550gat);
  nor x1676(s4607gat,s4554gat,s4551gat);
  nor x1677(s4611gat,s4491gat,s4557gat);
  nor x1678(s4612gat,s4557gat,s4488gat);
  nor x1679(s4613gat,s4561gat,s4562gat);
  nor x1680(s4616gat,s4563gat,s960gat);
  nor x1681(s4620gat,s4500gat,s4566gat);
  nor x1682(s4621gat,s4566gat,s1008gat);
  nor x1683(s4622gat,s4380gat,s4566gat);
  nor x1684(s4625gat,s4570gat,s4571gat);
  nor x1685(s4628gat,s4575gat,s4572gat);
  nor x1686(s4632gat,s4512gat,s4578gat);
  nor x1687(s4633gat,s4578gat,s4509gat);
  nor x1688(s4634gat,s4582gat,s4583gat);
  nor x1689(s4637gat,s4584gat,s1203gat);
  nor x1690(s4641gat,s4521gat,s4587gat);
  nor x1691(s4642gat,s4587gat,s1251gat);
  nor x1692(s4643gat,s4401gat,s4587gat);
  nor x1693(s4646gat,s4592gat,s4526gat);
  nor x1694(s4650gat,s4595gat,s4531gat);
  nor x1695(s4654gat,s4598gat,s4536gat);
  nor x1696(s4658gat,s4601gat,s4541gat);
  nor x1697(s4662gat,s4604gat,s4546gat);
  nor x1698(s4666gat,s4554gat,s4607gat);
  nor x1699(s4667gat,s4607gat,s4551gat);
  nor x1700(s4668gat,s4611gat,s4612gat);
  nor x1701(s4671gat,s4613gat,s912gat);
  nor x1702(s4675gat,s4563gat,s4616gat);
  nor x1703(s4676gat,s4616gat,s960gat);
  nor x1704(s4677gat,s4435gat,s4616gat);
  nor x1705(s4680gat,s4620gat,s4621gat);
  nor x1706(s4683gat,s4625gat,s4622gat);
  nor x1707(s4687gat,s4575gat,s4628gat);
  nor x1708(s4688gat,s4628gat,s4572gat);
  nor x1709(s4689gat,s4632gat,s4633gat);
  nor x1710(s4692gat,s4634gat,s1155gat);
  nor x1711(s4696gat,s4584gat,s4637gat);
  nor x1712(s4697gat,s4637gat,s1203gat);
  nor x1713(s4698gat,s4456gat,s4637gat);
  nor x1714(s4701gat,s4641gat,s4642gat);
  nor x1715(s4704gat,s1299gat,s4643gat);
  nor x1716(s4708gat,s4592gat,s4646gat);
  nor x1717(s4709gat,s4646gat,s4526gat);
  nor x1718(s4710gat,s4595gat,s4650gat);
  nor x1719(s4711gat,s4650gat,s4531gat);
  nor x1720(s4712gat,s4598gat,s4654gat);
  nor x1721(s4713gat,s4654gat,s4536gat);
  nor x1722(s4714gat,s4601gat,s4658gat);
  nor x1723(s4715gat,s4658gat,s4541gat);
  nor x1724(s4716gat,s4604gat,s4662gat);
  nor x1725(s4717gat,s4662gat,s4546gat);
  nor x1726(s4718gat,s4666gat,s4667gat);
  nor x1727(s4721gat,s4668gat,s864gat);
  nor x1728(s4725gat,s4613gat,s4671gat);
  nor x1729(s4726gat,s4671gat,s912gat);
  nor x1730(s4727gat,s4494gat,s4671gat);
  nor x1731(s4730gat,s4675gat,s4676gat);
  nor x1732(s4733gat,s4680gat,s4677gat);
  nor x1733(s4737gat,s4625gat,s4683gat);
  nor x1734(s4738gat,s4683gat,s4622gat);
  nor x1735(s4739gat,s4687gat,s4688gat);
  nor x1736(s4742gat,s4689gat,s1107gat);
  nor x1737(s4746gat,s4634gat,s4692gat);
  nor x1738(s4747gat,s4692gat,s1155gat);
  nor x1739(s4748gat,s4515gat,s4692gat);
  nor x1740(s4751gat,s4696gat,s4697gat);
  nor x1741(s4754gat,s4701gat,s4698gat);
  nor x1742(s4758gat,s1299gat,s4704gat);
  nor x1743(s4759gat,s4704gat,s4643gat);
  nor x1744(s4760gat,s4708gat,s4709gat);
  nor x1745(s4763gat,s4710gat,s4711gat);
  nor x1746(s4766gat,s4712gat,s4713gat);
  nor x1747(s4769gat,s4714gat,s4715gat);
  nor x1748(s4772gat,s4716gat,s4717gat);
  nor x1749(s4775gat,s4718gat,s816gat);
  nor x1750(s4779gat,s4668gat,s4721gat);
  nor x1751(s4780gat,s4721gat,s864gat);
  nor x1752(s4781gat,s4557gat,s4721gat);
  nor x1753(s4784gat,s4725gat,s4726gat);
  nor x1754(s4787gat,s4730gat,s4727gat);
  nor x1755(s4791gat,s4680gat,s4733gat);
  nor x1756(s4792gat,s4733gat,s4677gat);
  nor x1757(s4793gat,s4737gat,s4738gat);
  nor x1758(s4796gat,s4739gat,s1059gat);
  nor x1759(s4800gat,s4689gat,s4742gat);
  nor x1760(s4801gat,s4742gat,s1107gat);
  nor x1761(s4802gat,s4578gat,s4742gat);
  nor x1762(s4805gat,s4746gat,s4747gat);
  nor x1763(s4808gat,s4751gat,s4748gat);
  nor x1764(s4812gat,s4701gat,s4754gat);
  nor x1765(s4813gat,s4754gat,s4698gat);
  nor x1766(s4814gat,s4758gat,s4759gat);
  nor x1767(s4817gat,s4760gat,s576gat);
  nor x1768(s4821gat,s4763gat,s624gat);
  nor x1769(s4825gat,s4766gat,s672gat);
  nor x1770(s4829gat,s4769gat,s720gat);
  nor x1771(s4833gat,s4772gat,s768gat);
  nor x1772(s4837gat,s4718gat,s4775gat);
  nor x1773(s4838gat,s4775gat,s816gat);
  nor x1774(s4839gat,s4607gat,s4775gat);
  nor x1775(s4842gat,s4779gat,s4780gat);
  nor x1776(s4845gat,s4784gat,s4781gat);
  nor x1777(s4849gat,s4730gat,s4787gat);
  nor x1778(s4850gat,s4787gat,s4727gat);
  nor x1779(s4851gat,s4791gat,s4792gat);
  nor x1780(s4854gat,s4793gat,s1011gat);
  nor x1781(s4858gat,s4739gat,s4796gat);
  nor x1782(s4859gat,s4796gat,s1059gat);
  nor x1783(s4860gat,s4628gat,s4796gat);
  nor x1784(s4863gat,s4800gat,s4801gat);
  nor x1785(s4866gat,s4805gat,s4802gat);
  nor x1786(s4870gat,s4751gat,s4808gat);
  nor x1787(s4871gat,s4808gat,s4748gat);
  nor x1788(s4872gat,s4812gat,s4813gat);
  nor x1789(s4875gat,s4814gat,s1254gat);
  nor x1790(s4879gat,s4760gat,s4817gat);
  nor x1791(s4880gat,s4817gat,s576gat);
  nor x1792(s4881gat,s4646gat,s4817gat);
  nor x1793(s4884gat,s4763gat,s4821gat);
  nor x1794(s4885gat,s4821gat,s624gat);
  nor x1795(s4886gat,s4650gat,s4821gat);
  nor x1796(s4889gat,s4766gat,s4825gat);
  nor x1797(s4890gat,s4825gat,s672gat);
  nor x1798(s4891gat,s4654gat,s4825gat);
  nor x1799(s4894gat,s4769gat,s4829gat);
  nor x1800(s4895gat,s4829gat,s720gat);
  nor x1801(s4896gat,s4658gat,s4829gat);
  nor x1802(s4899gat,s4772gat,s4833gat);
  nor x1803(s4900gat,s4833gat,s768gat);
  nor x1804(s4901gat,s4662gat,s4833gat);
  nor x1805(s4904gat,s4837gat,s4838gat);
  nor x1806(s4907gat,s4842gat,s4839gat);
  nor x1807(s4911gat,s4784gat,s4845gat);
  nor x1808(s4912gat,s4845gat,s4781gat);
  nor x1809(s4913gat,s4849gat,s4850gat);
  nor x1810(s4916gat,s4851gat,s963gat);
  nor x1811(s4920gat,s4793gat,s4854gat);
  nor x1812(s4921gat,s4854gat,s1011gat);
  nor x1813(s4922gat,s4683gat,s4854gat);
  nor x1814(s4925gat,s4858gat,s4859gat);
  nor x1815(s4928gat,s4863gat,s4860gat);
  nor x1816(s4932gat,s4805gat,s4866gat);
  nor x1817(s4933gat,s4866gat,s4802gat);
  nor x1818(s4934gat,s4870gat,s4871gat);
  nor x1819(s4937gat,s4872gat,s1206gat);
  nor x1820(s4941gat,s4814gat,s4875gat);
  nor x1821(s4942gat,s4875gat,s1254gat);
  nor x1822(s4943gat,s4704gat,s4875gat);
  nor x1823(s4946gat,s4879gat,s4880gat);
  nor x1824(s4947gat,s4884gat,s4885gat);
  nor x1825(s4950gat,s4889gat,s4890gat);
  nor x1826(s4953gat,s4894gat,s4895gat);
  nor x1827(s4956gat,s4899gat,s4900gat);
  nor x1828(s4959gat,s4904gat,s4901gat);
  nor x1829(s4963gat,s4842gat,s4907gat);
  nor x1830(s4964gat,s4907gat,s4839gat);
  nor x1831(s4965gat,s4911gat,s4912gat);
  nor x1832(s4968gat,s4913gat,s915gat);
  nor x1833(s4972gat,s4851gat,s4916gat);
  nor x1834(s4973gat,s4916gat,s963gat);
  nor x1835(s4974gat,s4733gat,s4916gat);
  nor x1836(s4977gat,s4920gat,s4921gat);
  nor x1837(s4980gat,s4925gat,s4922gat);
  nor x1838(s4984gat,s4863gat,s4928gat);
  nor x1839(s4985gat,s4928gat,s4860gat);
  nor x1840(s4986gat,s4932gat,s4933gat);
  nor x1841(s4989gat,s4934gat,s1158gat);
  nor x1842(s4993gat,s4872gat,s4937gat);
  nor x1843(s4994gat,s4937gat,s1206gat);
  nor x1844(s4995gat,s4754gat,s4937gat);
  nor x1845(s4998gat,s4941gat,s4942gat);
  nor x1846(s5001gat,s1302gat,s4943gat);
  nor x1847(s5005gat,s4947gat,s4881gat);
  nor x1848(s5009gat,s4950gat,s4886gat);
  nor x1849(s5013gat,s4953gat,s4891gat);
  nor x1850(s5017gat,s4956gat,s4896gat);
  nor x1851(s5021gat,s4904gat,s4959gat);
  nor x1852(s5022gat,s4959gat,s4901gat);
  nor x1853(s5023gat,s4963gat,s4964gat);
  nor x1854(s5026gat,s4965gat,s867gat);
  nor x1855(s5030gat,s4913gat,s4968gat);
  nor x1856(s5031gat,s4968gat,s915gat);
  nor x1857(s5032gat,s4787gat,s4968gat);
  nor x1858(s5035gat,s4972gat,s4973gat);
  nor x1859(s5038gat,s4977gat,s4974gat);
  nor x1860(s5042gat,s4925gat,s4980gat);
  nor x1861(s5043gat,s4980gat,s4922gat);
  nor x1862(s5044gat,s4984gat,s4985gat);
  nor x1863(s5047gat,s4986gat,s1110gat);
  nor x1864(s5051gat,s4934gat,s4989gat);
  nor x1865(s5052gat,s4989gat,s1158gat);
  nor x1866(s5053gat,s4808gat,s4989gat);
  nor x1867(s5056gat,s4993gat,s4994gat);
  nor x1868(s5059gat,s4998gat,s4995gat);
  nor x1869(s5063gat,s1302gat,s5001gat);
  nor x1870(s5064gat,s5001gat,s4943gat);
  nor x1871(s5065gat,s4947gat,s5005gat);
  nor x1872(s5066gat,s5005gat,s4881gat);
  nor x1873(s5067gat,s4950gat,s5009gat);
  nor x1874(s5068gat,s5009gat,s4886gat);
  nor x1875(s5069gat,s4953gat,s5013gat);
  nor x1876(s5070gat,s5013gat,s4891gat);
  nor x1877(s5071gat,s4956gat,s5017gat);
  nor x1878(s5072gat,s5017gat,s4896gat);
  nor x1879(s5073gat,s5021gat,s5022gat);
  nor x1880(s5076gat,s5023gat,s819gat);
  nor x1881(s5080gat,s4965gat,s5026gat);
  nor x1882(s5081gat,s5026gat,s867gat);
  nor x1883(s5082gat,s4845gat,s5026gat);
  nor x1884(s5085gat,s5030gat,s5031gat);
  nor x1885(s5088gat,s5035gat,s5032gat);
  nor x1886(s5092gat,s4977gat,s5038gat);
  nor x1887(s5093gat,s5038gat,s4974gat);
  nor x1888(s5094gat,s5042gat,s5043gat);
  nor x1889(s5097gat,s5044gat,s1062gat);
  nor x1890(s5101gat,s4986gat,s5047gat);
  nor x1891(s5102gat,s5047gat,s1110gat);
  nor x1892(s5103gat,s4866gat,s5047gat);
  nor x1893(s5106gat,s5051gat,s5052gat);
  nor x1894(s5109gat,s5056gat,s5053gat);
  nor x1895(s5113gat,s4998gat,s5059gat);
  nor x1896(s5114gat,s5059gat,s4995gat);
  nor x1897(s5115gat,s5063gat,s5064gat);
  nor x1898(s5118gat,s5065gat,s5066gat);
  nor x1899(s5121gat,s5067gat,s5068gat);
  nor x1900(s5124gat,s5069gat,s5070gat);
  nor x1901(s5127gat,s5071gat,s5072gat);
  nor x1902(s5130gat,s5073gat,s771gat);
  nor x1903(s5134gat,s5023gat,s5076gat);
  nor x1904(s5135gat,s5076gat,s819gat);
  nor x1905(s5136gat,s4907gat,s5076gat);
  nor x1906(s5139gat,s5080gat,s5081gat);
  nor x1907(s5142gat,s5085gat,s5082gat);
  nor x1908(s5146gat,s5035gat,s5088gat);
  nor x1909(s5147gat,s5088gat,s5032gat);
  nor x1910(s5148gat,s5092gat,s5093gat);
  nor x1911(s5151gat,s5094gat,s1014gat);
  nor x1912(s5155gat,s5044gat,s5097gat);
  nor x1913(s5156gat,s5097gat,s1062gat);
  nor x1914(s5157gat,s4928gat,s5097gat);
  nor x1915(s5160gat,s5101gat,s5102gat);
  nor x1916(s5163gat,s5106gat,s5103gat);
  nor x1917(s5167gat,s5056gat,s5109gat);
  nor x1918(s5168gat,s5109gat,s5053gat);
  nor x1919(s5169gat,s5113gat,s5114gat);
  nor x1920(s5172gat,s5115gat,s1257gat);
  nor x1921(s5176gat,s5118gat,s579gat);
  nor x1922(s5180gat,s5121gat,s627gat);
  nor x1923(s5184gat,s5124gat,s675gat);
  nor x1924(s5188gat,s5127gat,s723gat);
  nor x1925(s5192gat,s5073gat,s5130gat);
  nor x1926(s5193gat,s5130gat,s771gat);
  nor x1927(s5194gat,s4959gat,s5130gat);
  nor x1928(s5197gat,s5134gat,s5135gat);
  nor x1929(s5200gat,s5139gat,s5136gat);
  nor x1930(s5204gat,s5085gat,s5142gat);
  nor x1931(s5205gat,s5142gat,s5082gat);
  nor x1932(s5206gat,s5146gat,s5147gat);
  nor x1933(s5209gat,s5148gat,s966gat);
  nor x1934(s5213gat,s5094gat,s5151gat);
  nor x1935(s5214gat,s5151gat,s1014gat);
  nor x1936(s5215gat,s4980gat,s5151gat);
  nor x1937(s5218gat,s5155gat,s5156gat);
  nor x1938(s5221gat,s5160gat,s5157gat);
  nor x1939(s5225gat,s5106gat,s5163gat);
  nor x1940(s5226gat,s5163gat,s5103gat);
  nor x1941(s5227gat,s5167gat,s5168gat);
  nor x1942(s5230gat,s5169gat,s1209gat);
  nor x1943(s5234gat,s5115gat,s5172gat);
  nor x1944(s5235gat,s5172gat,s1257gat);
  nor x1945(s5236gat,s5001gat,s5172gat);
  nor x1946(s5239gat,s5118gat,s5176gat);
  nor x1947(s5240gat,s5176gat,s579gat);
  nor x1948(s5241gat,s5005gat,s5176gat);
  nor x1949(s5244gat,s5121gat,s5180gat);
  nor x1950(s5245gat,s5180gat,s627gat);
  nor x1951(s5246gat,s5009gat,s5180gat);
  nor x1952(s5249gat,s5124gat,s5184gat);
  nor x1953(s5250gat,s5184gat,s675gat);
  nor x1954(s5251gat,s5013gat,s5184gat);
  nor x1955(s5254gat,s5127gat,s5188gat);
  nor x1956(s5255gat,s5188gat,s723gat);
  nor x1957(s5256gat,s5017gat,s5188gat);
  nor x1958(s5259gat,s5192gat,s5193gat);
  nor x1959(s5262gat,s5197gat,s5194gat);
  nor x1960(s5266gat,s5139gat,s5200gat);
  nor x1961(s5267gat,s5200gat,s5136gat);
  nor x1962(s5268gat,s5204gat,s5205gat);
  nor x1963(s5271gat,s5206gat,s918gat);
  nor x1964(s5275gat,s5148gat,s5209gat);
  nor x1965(s5276gat,s5209gat,s966gat);
  nor x1966(s5277gat,s5038gat,s5209gat);
  nor x1967(s5280gat,s5213gat,s5214gat);
  nor x1968(s5283gat,s5218gat,s5215gat);
  nor x1969(s5287gat,s5160gat,s5221gat);
  nor x1970(s5288gat,s5221gat,s5157gat);
  nor x1971(s5289gat,s5225gat,s5226gat);
  nor x1972(s5292gat,s5227gat,s1161gat);
  nor x1973(s5296gat,s5169gat,s5230gat);
  nor x1974(s5297gat,s5230gat,s1209gat);
  nor x1975(s5298gat,s5059gat,s5230gat);
  nor x1976(s5301gat,s5234gat,s5235gat);
  nor x1977(s5304gat,s1305gat,s5236gat);
  nor x1978(s5308gat,s5239gat,s5240gat);
  nor x1979(s5309gat,s5244gat,s5245gat);
  nor x1980(s5312gat,s5249gat,s5250gat);
  nor x1981(s5315gat,s5254gat,s5255gat);
  nor x1982(s5318gat,s5259gat,s5256gat);
  nor x1983(s5322gat,s5197gat,s5262gat);
  nor x1984(s5323gat,s5262gat,s5194gat);
  nor x1985(s5324gat,s5266gat,s5267gat);
  nor x1986(s5327gat,s5268gat,s870gat);
  nor x1987(s5331gat,s5206gat,s5271gat);
  nor x1988(s5332gat,s5271gat,s918gat);
  nor x1989(s5333gat,s5088gat,s5271gat);
  nor x1990(s5336gat,s5275gat,s5276gat);
  nor x1991(s5339gat,s5280gat,s5277gat);
  nor x1992(s5343gat,s5218gat,s5283gat);
  nor x1993(s5344gat,s5283gat,s5215gat);
  nor x1994(s5345gat,s5287gat,s5288gat);
  nor x1995(s5348gat,s5289gat,s1113gat);
  nor x1996(s5352gat,s5227gat,s5292gat);
  nor x1997(s5353gat,s5292gat,s1161gat);
  nor x1998(s5354gat,s5109gat,s5292gat);
  nor x1999(s5357gat,s5296gat,s5297gat);
  nor x2000(s5360gat,s5301gat,s5298gat);
  nor x2001(s5364gat,s1305gat,s5304gat);
  nor x2002(s5365gat,s5304gat,s5236gat);
  nor x2003(s5366gat,s5309gat,s5241gat);
  nor x2004(s5370gat,s5312gat,s5246gat);
  nor x2005(s5374gat,s5315gat,s5251gat);
  nor x2006(s5378gat,s5259gat,s5318gat);
  nor x2007(s5379gat,s5318gat,s5256gat);
  nor x2008(s5380gat,s5322gat,s5323gat);
  nor x2009(s5383gat,s5324gat,s822gat);
  nor x2010(s5387gat,s5268gat,s5327gat);
  nor x2011(s5388gat,s5327gat,s870gat);
  nor x2012(s5389gat,s5142gat,s5327gat);
  nor x2013(s5392gat,s5331gat,s5332gat);
  nor x2014(s5395gat,s5336gat,s5333gat);
  nor x2015(s5399gat,s5280gat,s5339gat);
  nor x2016(s5400gat,s5339gat,s5277gat);
  nor x2017(s5401gat,s5343gat,s5344gat);
  nor x2018(s5404gat,s5345gat,s1065gat);
  nor x2019(s5408gat,s5289gat,s5348gat);
  nor x2020(s5409gat,s5348gat,s1113gat);
  nor x2021(s5410gat,s5163gat,s5348gat);
  nor x2022(s5413gat,s5352gat,s5353gat);
  nor x2023(s5416gat,s5357gat,s5354gat);
  nor x2024(s5420gat,s5301gat,s5360gat);
  nor x2025(s5421gat,s5360gat,s5298gat);
  nor x2026(s5422gat,s5364gat,s5365gat);
  nor x2027(s5425gat,s5309gat,s5366gat);
  nor x2028(s5426gat,s5366gat,s5241gat);
  nor x2029(s5427gat,s5312gat,s5370gat);
  nor x2030(s5428gat,s5370gat,s5246gat);
  nor x2031(s5429gat,s5315gat,s5374gat);
  nor x2032(s5430gat,s5374gat,s5251gat);
  nor x2033(s5431gat,s5378gat,s5379gat);
  nor x2034(s5434gat,s5380gat,s774gat);
  nor x2035(s5438gat,s5324gat,s5383gat);
  nor x2036(s5439gat,s5383gat,s822gat);
  nor x2037(s5440gat,s5200gat,s5383gat);
  nor x2038(s5443gat,s5387gat,s5388gat);
  nor x2039(s5446gat,s5392gat,s5389gat);
  nor x2040(s5450gat,s5336gat,s5395gat);
  nor x2041(s5451gat,s5395gat,s5333gat);
  nor x2042(s5452gat,s5399gat,s5400gat);
  nor x2043(s5455gat,s5401gat,s1017gat);
  nor x2044(s5459gat,s5345gat,s5404gat);
  nor x2045(s5460gat,s5404gat,s1065gat);
  nor x2046(s5461gat,s5221gat,s5404gat);
  nor x2047(s5464gat,s5408gat,s5409gat);
  nor x2048(s5467gat,s5413gat,s5410gat);
  nor x2049(s5471gat,s5357gat,s5416gat);
  nor x2050(s5472gat,s5416gat,s5354gat);
  nor x2051(s5473gat,s5420gat,s5421gat);
  nor x2052(s5476gat,s5422gat,s1260gat);
  nor x2053(s5480gat,s5425gat,s5426gat);
  nor x2054(s5483gat,s5427gat,s5428gat);
  nor x2055(s5486gat,s5429gat,s5430gat);
  nor x2056(s5489gat,s5431gat,s726gat);
  nor x2057(s5493gat,s5380gat,s5434gat);
  nor x2058(s5494gat,s5434gat,s774gat);
  nor x2059(s5495gat,s5262gat,s5434gat);
  nor x2060(s5498gat,s5438gat,s5439gat);
  nor x2061(s5501gat,s5443gat,s5440gat);
  nor x2062(s5505gat,s5392gat,s5446gat);
  nor x2063(s5506gat,s5446gat,s5389gat);
  nor x2064(s5507gat,s5450gat,s5451gat);
  nor x2065(s5510gat,s5452gat,s969gat);
  nor x2066(s5514gat,s5401gat,s5455gat);
  nor x2067(s5515gat,s5455gat,s1017gat);
  nor x2068(s5516gat,s5283gat,s5455gat);
  nor x2069(s5519gat,s5459gat,s5460gat);
  nor x2070(s5522gat,s5464gat,s5461gat);
  nor x2071(s5526gat,s5413gat,s5467gat);
  nor x2072(s5527gat,s5467gat,s5410gat);
  nor x2073(s5528gat,s5471gat,s5472gat);
  nor x2074(s5531gat,s5473gat,s1212gat);
  nor x2075(s5535gat,s5422gat,s5476gat);
  nor x2076(s5536gat,s5476gat,s1260gat);
  nor x2077(s5537gat,s5304gat,s5476gat);
  nor x2078(s5540gat,s5480gat,s582gat);
  nor x2079(s5544gat,s5483gat,s630gat);
  nor x2080(s5548gat,s5486gat,s678gat);
  nor x2081(s5552gat,s5431gat,s5489gat);
  nor x2082(s5553gat,s5489gat,s726gat);
  nor x2083(s5554gat,s5318gat,s5489gat);
  nor x2084(s5557gat,s5493gat,s5494gat);
  nor x2085(s5560gat,s5498gat,s5495gat);
  nor x2086(s5564gat,s5443gat,s5501gat);
  nor x2087(s5565gat,s5501gat,s5440gat);
  nor x2088(s5566gat,s5505gat,s5506gat);
  nor x2089(s5569gat,s5507gat,s921gat);
  nor x2090(s5573gat,s5452gat,s5510gat);
  nor x2091(s5574gat,s5510gat,s969gat);
  nor x2092(s5575gat,s5339gat,s5510gat);
  nor x2093(s5578gat,s5514gat,s5515gat);
  nor x2094(s5581gat,s5519gat,s5516gat);
  nor x2095(s5585gat,s5464gat,s5522gat);
  nor x2096(s5586gat,s5522gat,s5461gat);
  nor x2097(s5587gat,s5526gat,s5527gat);
  nor x2098(s5590gat,s5528gat,s1164gat);
  nor x2099(s5594gat,s5473gat,s5531gat);
  nor x2100(s5595gat,s5531gat,s1212gat);
  nor x2101(s5596gat,s5360gat,s5531gat);
  nor x2102(s5599gat,s5535gat,s5536gat);
  nor x2103(s5602gat,s1308gat,s5537gat);
  nor x2104(s5606gat,s5480gat,s5540gat);
  nor x2105(s5607gat,s5540gat,s582gat);
  nor x2106(s5608gat,s5366gat,s5540gat);
  nor x2107(s5611gat,s5483gat,s5544gat);
  nor x2108(s5612gat,s5544gat,s630gat);
  nor x2109(s5613gat,s5370gat,s5544gat);
  nor x2110(s5616gat,s5486gat,s5548gat);
  nor x2111(s5617gat,s5548gat,s678gat);
  nor x2112(s5618gat,s5374gat,s5548gat);
  nor x2113(s5621gat,s5552gat,s5553gat);
  nor x2114(s5624gat,s5557gat,s5554gat);
  nor x2115(s5628gat,s5498gat,s5560gat);
  nor x2116(s5629gat,s5560gat,s5495gat);
  nor x2117(s5630gat,s5564gat,s5565gat);
  nor x2118(s5633gat,s5566gat,s873gat);
  nor x2119(s5637gat,s5507gat,s5569gat);
  nor x2120(s5638gat,s5569gat,s921gat);
  nor x2121(s5639gat,s5395gat,s5569gat);
  nor x2122(s5642gat,s5573gat,s5574gat);
  nor x2123(s5645gat,s5578gat,s5575gat);
  nor x2124(s5649gat,s5519gat,s5581gat);
  nor x2125(s5650gat,s5581gat,s5516gat);
  nor x2126(s5651gat,s5585gat,s5586gat);
  nor x2127(s5654gat,s5587gat,s1116gat);
  nor x2128(s5658gat,s5528gat,s5590gat);
  nor x2129(s5659gat,s5590gat,s1164gat);
  nor x2130(s5660gat,s5416gat,s5590gat);
  nor x2131(s5663gat,s5594gat,s5595gat);
  nor x2132(s5666gat,s5599gat,s5596gat);
  nor x2133(s5670gat,s1308gat,s5602gat);
  nor x2134(s5671gat,s5602gat,s5537gat);
  nor x2135(s5672gat,s5606gat,s5607gat);
  nor x2136(s5673gat,s5611gat,s5612gat);
  nor x2137(s5676gat,s5616gat,s5617gat);
  nor x2138(s5679gat,s5621gat,s5618gat);
  nor x2139(s5683gat,s5557gat,s5624gat);
  nor x2140(s5684gat,s5624gat,s5554gat);
  nor x2141(s5685gat,s5628gat,s5629gat);
  nor x2142(s5688gat,s5630gat,s825gat);
  nor x2143(s5692gat,s5566gat,s5633gat);
  nor x2144(s5693gat,s5633gat,s873gat);
  nor x2145(s5694gat,s5446gat,s5633gat);
  nor x2146(s5697gat,s5637gat,s5638gat);
  nor x2147(s5700gat,s5642gat,s5639gat);
  nor x2148(s5704gat,s5578gat,s5645gat);
  nor x2149(s5705gat,s5645gat,s5575gat);
  nor x2150(s5706gat,s5649gat,s5650gat);
  nor x2151(s5709gat,s5651gat,s1068gat);
  nor x2152(s5713gat,s5587gat,s5654gat);
  nor x2153(s5714gat,s5654gat,s1116gat);
  nor x2154(s5715gat,s5467gat,s5654gat);
  nor x2155(s5718gat,s5658gat,s5659gat);
  nor x2156(s5721gat,s5663gat,s5660gat);
  nor x2157(s5725gat,s5599gat,s5666gat);
  nor x2158(s5726gat,s5666gat,s5596gat);
  nor x2159(s5727gat,s5670gat,s5671gat);
  nor x2160(s5730gat,s5673gat,s5608gat);
  nor x2161(s5734gat,s5676gat,s5613gat);
  nor x2162(s5738gat,s5621gat,s5679gat);
  nor x2163(s5739gat,s5679gat,s5618gat);
  nor x2164(s5740gat,s5683gat,s5684gat);
  nor x2165(s5743gat,s5685gat,s777gat);
  nor x2166(s5747gat,s5630gat,s5688gat);
  nor x2167(s5748gat,s5688gat,s825gat);
  nor x2168(s5749gat,s5501gat,s5688gat);
  nor x2169(s5752gat,s5692gat,s5693gat);
  nor x2170(s5755gat,s5697gat,s5694gat);
  nor x2171(s5759gat,s5642gat,s5700gat);
  nor x2172(s5760gat,s5700gat,s5639gat);
  nor x2173(s5761gat,s5704gat,s5705gat);
  nor x2174(s5764gat,s5706gat,s1020gat);
  nor x2175(s5768gat,s5651gat,s5709gat);
  nor x2176(s5769gat,s5709gat,s1068gat);
  nor x2177(s5770gat,s5522gat,s5709gat);
  nor x2178(s5773gat,s5713gat,s5714gat);
  nor x2179(s5776gat,s5718gat,s5715gat);
  nor x2180(s5780gat,s5663gat,s5721gat);
  nor x2181(s5781gat,s5721gat,s5660gat);
  nor x2182(s5782gat,s5725gat,s5726gat);
  nor x2183(s5785gat,s5673gat,s5730gat);
  nor x2184(s5786gat,s5730gat,s5608gat);
  nor x2185(s5787gat,s5676gat,s5734gat);
  nor x2186(s5788gat,s5734gat,s5613gat);
  nor x2187(s5789gat,s5738gat,s5739gat);
  nor x2188(s5792gat,s5740gat,s729gat);
  nor x2189(s5796gat,s5685gat,s5743gat);
  nor x2190(s5797gat,s5743gat,s777gat);
  nor x2191(s5798gat,s5560gat,s5743gat);
  nor x2192(s5801gat,s5747gat,s5748gat);
  nor x2193(s5804gat,s5752gat,s5749gat);
  nor x2194(s5808gat,s5697gat,s5755gat);
  nor x2195(s5809gat,s5755gat,s5694gat);
  nor x2196(s5810gat,s5759gat,s5760gat);
  nor x2197(s5813gat,s5761gat,s972gat);
  nor x2198(s5817gat,s5706gat,s5764gat);
  nor x2199(s5818gat,s5764gat,s1020gat);
  nor x2200(s5819gat,s5581gat,s5764gat);
  nor x2201(s5822gat,s5768gat,s5769gat);
  nor x2202(s5825gat,s5773gat,s5770gat);
  nor x2203(s5829gat,s5718gat,s5776gat);
  nor x2204(s5830gat,s5776gat,s5715gat);
  nor x2205(s5831gat,s5780gat,s5781gat);
  nor x2206(s5834gat,s5785gat,s5786gat);
  nor x2207(s5837gat,s5787gat,s5788gat);
  nor x2208(s5840gat,s5789gat,s681gat);
  nor x2209(s5844gat,s5740gat,s5792gat);
  nor x2210(s5845gat,s5792gat,s729gat);
  nor x2211(s5846gat,s5624gat,s5792gat);
  nor x2212(s5849gat,s5796gat,s5797gat);
  nor x2213(s5852gat,s5801gat,s5798gat);
  nor x2214(s5856gat,s5752gat,s5804gat);
  nor x2215(s5857gat,s5804gat,s5749gat);
  nor x2216(s5858gat,s5808gat,s5809gat);
  nor x2217(s5861gat,s5810gat,s924gat);
  nor x2218(s5865gat,s5761gat,s5813gat);
  nor x2219(s5866gat,s5813gat,s972gat);
  nor x2220(s5867gat,s5645gat,s5813gat);
  nor x2221(s5870gat,s5817gat,s5818gat);
  nor x2222(s5873gat,s5822gat,s5819gat);
  nor x2223(s5877gat,s5773gat,s5825gat);
  nor x2224(s5878gat,s5825gat,s5770gat);
  nor x2225(s5879gat,s5829gat,s5830gat);
  nor x2226(s5882gat,s5834gat,s585gat);
  nor x2227(s5886gat,s5837gat,s633gat);
  nor x2228(s5890gat,s5789gat,s5840gat);
  nor x2229(s5891gat,s5840gat,s681gat);
  nor x2230(s5892gat,s5679gat,s5840gat);
  nor x2231(s5895gat,s5844gat,s5845gat);
  nor x2232(s5898gat,s5849gat,s5846gat);
  nor x2233(s5902gat,s5801gat,s5852gat);
  nor x2234(s5903gat,s5852gat,s5798gat);
  nor x2235(s5904gat,s5856gat,s5857gat);
  nor x2236(s5907gat,s5858gat,s876gat);
  nor x2237(s5911gat,s5810gat,s5861gat);
  nor x2238(s5912gat,s5861gat,s924gat);
  nor x2239(s5913gat,s5700gat,s5861gat);
  nor x2240(s5916gat,s5865gat,s5866gat);
  nor x2241(s5919gat,s5870gat,s5867gat);
  nor x2242(s5923gat,s5822gat,s5873gat);
  nor x2243(s5924gat,s5873gat,s5819gat);
  nor x2244(s5925gat,s5877gat,s5878gat);
  nor x2245(s5928gat,s5834gat,s5882gat);
  nor x2246(s5929gat,s5882gat,s585gat);
  nor x2247(s5930gat,s5730gat,s5882gat);
  nor x2248(s5933gat,s5837gat,s5886gat);
  nor x2249(s5934gat,s5886gat,s633gat);
  nor x2250(s5935gat,s5734gat,s5886gat);
  nor x2251(s5938gat,s5890gat,s5891gat);
  nor x2252(s5941gat,s5895gat,s5892gat);
  nor x2253(s5945gat,s5849gat,s5898gat);
  nor x2254(s5946gat,s5898gat,s5846gat);
  nor x2255(s5947gat,s5902gat,s5903gat);
  nor x2256(s5950gat,s5904gat,s828gat);
  nor x2257(s5954gat,s5858gat,s5907gat);
  nor x2258(s5955gat,s5907gat,s876gat);
  nor x2259(s5956gat,s5755gat,s5907gat);
  nor x2260(s5959gat,s5911gat,s5912gat);
  nor x2261(s5962gat,s5916gat,s5913gat);
  nor x2262(s5966gat,s5870gat,s5919gat);
  nor x2263(s5967gat,s5919gat,s5867gat);
  nor x2264(s5968gat,s5923gat,s5924gat);
  nor x2265(s5971gat,s5928gat,s5929gat);
  nor x2266(s5972gat,s5933gat,s5934gat);
  nor x2267(s5975gat,s5938gat,s5935gat);
  nor x2268(s5979gat,s5895gat,s5941gat);
  nor x2269(s5980gat,s5941gat,s5892gat);
  nor x2270(s5981gat,s5945gat,s5946gat);
  nor x2271(s5984gat,s5947gat,s780gat);
  nor x2272(s5988gat,s5904gat,s5950gat);
  nor x2273(s5989gat,s5950gat,s828gat);
  nor x2274(s5990gat,s5804gat,s5950gat);
  nor x2275(s5993gat,s5954gat,s5955gat);
  nor x2276(s5996gat,s5959gat,s5956gat);
  nor x2277(s6000gat,s5916gat,s5962gat);
  nor x2278(s6001gat,s5962gat,s5913gat);
  nor x2279(s6002gat,s5966gat,s5967gat);
  nor x2280(s6005gat,s5972gat,s5930gat);
  nor x2281(s6009gat,s5938gat,s5975gat);
  nor x2282(s6010gat,s5975gat,s5935gat);
  nor x2283(s6011gat,s5979gat,s5980gat);
  nor x2284(s6014gat,s5981gat,s732gat);
  nor x2285(s6018gat,s5947gat,s5984gat);
  nor x2286(s6019gat,s5984gat,s780gat);
  nor x2287(s6020gat,s5852gat,s5984gat);
  nor x2288(s6023gat,s5988gat,s5989gat);
  nor x2289(s6026gat,s5993gat,s5990gat);
  nor x2290(s6030gat,s5959gat,s5996gat);
  nor x2291(s6031gat,s5996gat,s5956gat);
  nor x2292(s6032gat,s6000gat,s6001gat);
  nor x2293(s6035gat,s5972gat,s6005gat);
  nor x2294(s6036gat,s6005gat,s5930gat);
  nor x2295(s6037gat,s6009gat,s6010gat);
  nor x2296(s6040gat,s6011gat,s684gat);
  nor x2297(s6044gat,s5981gat,s6014gat);
  nor x2298(s6045gat,s6014gat,s732gat);
  nor x2299(s6046gat,s5898gat,s6014gat);
  nor x2300(s6049gat,s6018gat,s6019gat);
  nor x2301(s6052gat,s6023gat,s6020gat);
  nor x2302(s6056gat,s5993gat,s6026gat);
  nor x2303(s6057gat,s6026gat,s5990gat);
  nor x2304(s6058gat,s6030gat,s6031gat);
  nor x2305(s6061gat,s6035gat,s6036gat);
  nor x2306(s6064gat,s6037gat,s636gat);
  nor x2307(s6068gat,s6011gat,s6040gat);
  nor x2308(s6069gat,s6040gat,s684gat);
  nor x2309(s6070gat,s5941gat,s6040gat);
  nor x2310(s6073gat,s6044gat,s6045gat);
  nor x2311(s6076gat,s6049gat,s6046gat);
  nor x2312(s6080gat,s6023gat,s6052gat);
  nor x2313(s6081gat,s6052gat,s6020gat);
  nor x2314(s6082gat,s6056gat,s6057gat);
  nor x2315(s6085gat,s6061gat,s588gat);
  nor x2316(s6089gat,s6037gat,s6064gat);
  nor x2317(s6090gat,s6064gat,s636gat);
  nor x2318(s6091gat,s5975gat,s6064gat);
  nor x2319(s6094gat,s6068gat,s6069gat);
  nor x2320(s6097gat,s6073gat,s6070gat);
  nor x2321(s6101gat,s6049gat,s6076gat);
  nor x2322(s6102gat,s6076gat,s6046gat);
  nor x2323(s6103gat,s6080gat,s6081gat);
  nor x2324(s6106gat,s6061gat,s6085gat);
  nor x2325(s6107gat,s6085gat,s588gat);
  nor x2326(s6108gat,s6005gat,s6085gat);
  nor x2327(s6111gat,s6089gat,s6090gat);
  nor x2328(s6114gat,s6094gat,s6091gat);
  nor x2329(s6118gat,s6073gat,s6097gat);
  nor x2330(s6119gat,s6097gat,s6070gat);
  nor x2331(s6120gat,s6101gat,s6102gat);
  nor x2332(s6123gat,s6106gat,s6107gat);
  nor x2333(s6124gat,s6111gat,s6108gat);
  nor x2334(s6128gat,s6094gat,s6114gat);
  nor x2335(s6129gat,s6114gat,s6091gat);
  nor x2336(s6130gat,s6118gat,s6119gat);
  nor x2337(s6133gat,s6111gat,s6124gat);
  nor x2338(s6134gat,s6124gat,s6108gat);
  nor x2339(s6135gat,s6128gat,s6129gat);
  nor x2340(s6138gat,s6133gat,s6134gat);
  not x2341(s6141gat,s6138gat);
  nor x2342(s6145gat,s6138gat,s6141gat);
  not x2343(s6146gat,s6141gat);
  nor x2344(s6147gat,s6124gat,s6141gat);
  nor x2345(s6150gat,s6145gat,s6146gat);
  nor x2346(s6151gat,s6135gat,s6147gat);
  nor x2347(s6155gat,s6135gat,s6151gat);
  nor x2348(s6156gat,s6151gat,s6147gat);
  nor x2349(s6157gat,s6114gat,s6151gat);
  nor x2350(s6160gat,s6155gat,s6156gat);
  nor x2351(s6161gat,s6130gat,s6157gat);
  nor x2352(s6165gat,s6130gat,s6161gat);
  nor x2353(s6166gat,s6161gat,s6157gat);
  nor x2354(s6167gat,s6097gat,s6161gat);
  nor x2355(s6170gat,s6165gat,s6166gat);
  nor x2356(s6171gat,s6120gat,s6167gat);
  nor x2357(s6175gat,s6120gat,s6171gat);
  nor x2358(s6176gat,s6171gat,s6167gat);
  nor x2359(s6177gat,s6076gat,s6171gat);
  nor x2360(s6180gat,s6175gat,s6176gat);
  nor x2361(s6181gat,s6103gat,s6177gat);
  nor x2362(s6185gat,s6103gat,s6181gat);
  nor x2363(s6186gat,s6181gat,s6177gat);
  nor x2364(s6187gat,s6052gat,s6181gat);
  nor x2365(s6190gat,s6185gat,s6186gat);
  nor x2366(s6191gat,s6082gat,s6187gat);
  nor x2367(s6195gat,s6082gat,s6191gat);
  nor x2368(s6196gat,s6191gat,s6187gat);
  nor x2369(s6197gat,s6026gat,s6191gat);
  nor x2370(s6200gat,s6195gat,s6196gat);
  nor x2371(s6201gat,s6058gat,s6197gat);
  nor x2372(s6205gat,s6058gat,s6201gat);
  nor x2373(s6206gat,s6201gat,s6197gat);
  nor x2374(s6207gat,s5996gat,s6201gat);
  nor x2375(s6210gat,s6205gat,s6206gat);
  nor x2376(s6211gat,s6032gat,s6207gat);
  nor x2377(s6215gat,s6032gat,s6211gat);
  nor x2378(s6216gat,s6211gat,s6207gat);
  nor x2379(s6217gat,s5962gat,s6211gat);
  nor x2380(s6220gat,s6215gat,s6216gat);
  nor x2381(s6221gat,s6002gat,s6217gat);
  nor x2382(s6225gat,s6002gat,s6221gat);
  nor x2383(s6226gat,s6221gat,s6217gat);
  nor x2384(s6227gat,s5919gat,s6221gat);
  nor x2385(s6230gat,s6225gat,s6226gat);
  nor x2386(s6231gat,s5968gat,s6227gat);
  nor x2387(s6235gat,s5968gat,s6231gat);
  nor x2388(s6236gat,s6231gat,s6227gat);
  nor x2389(s6237gat,s5873gat,s6231gat);
  nor x2390(s6240gat,s6235gat,s6236gat);
  nor x2391(s6241gat,s5925gat,s6237gat);
  nor x2392(s6245gat,s5925gat,s6241gat);
  nor x2393(s6246gat,s6241gat,s6237gat);
  nor x2394(s6247gat,s5825gat,s6241gat);
  nor x2395(s6250gat,s6245gat,s6246gat);
  nor x2396(s6251gat,s5879gat,s6247gat);
  nor x2397(s6255gat,s5879gat,s6251gat);
  nor x2398(s6256gat,s6251gat,s6247gat);
  nor x2399(s6257gat,s5776gat,s6251gat);
  nor x2400(s6260gat,s6255gat,s6256gat);
  nor x2401(s6261gat,s5831gat,s6257gat);
  nor x2402(s6265gat,s5831gat,s6261gat);
  nor x2403(s6266gat,s6261gat,s6257gat);
  nor x2404(s6267gat,s5721gat,s6261gat);
  nor x2405(s6270gat,s6265gat,s6266gat);
  nor x2406(s6271gat,s5782gat,s6267gat);
  nor x2407(s6275gat,s5782gat,s6271gat);
  nor x2408(s6276gat,s6271gat,s6267gat);
  nor x2409(s6277gat,s5666gat,s6271gat);
  nor x2410(s6280gat,s6275gat,s6276gat);
  nor x2411(s6281gat,s5727gat,s6277gat);
  nor x2412(s6285gat,s5727gat,s6281gat);
  nor x2413(s6286gat,s6281gat,s6277gat);
  nor x2414(s6287gat,s5602gat,s6281gat);
  nor x2415(s6288gat,s6285gat,s6286gat);

endmodule
